// soc_system.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module soc_system (
		input  wire [1:0]  button_pio_export,                     //                button_pio.export
		input  wire        clk_clk,                               //                       clk.clk
		input  wire [3:0]  dipsw_pio_export,                      //                 dipsw_pio.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,      //  hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,     // hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,  //   hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,      //  hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_clk_clk,                     //             hps_0_h2f_clk.clk
		output wire        hps_0_h2f_reset_reset_n,               //           hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, //              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //                          .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //                          .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //                          .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //                          .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //                          .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //                          .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //                          .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //                          .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //                          .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //                          .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //                          .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //                          .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //                          .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //                          .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //                          .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //                          .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //                          .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //                          .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //                          .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //                          .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //                          .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //                          .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //                          .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //                          .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //                          .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //                          .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //                          .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //                          .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //                          .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //                          .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //                          .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,    //                          .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,   //                          .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,   //                          .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,    //                          .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //                          .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //                          .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //                          .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //                          .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,     //                          .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,     //                          .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //                          .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //                          .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,  //                          .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  //                          .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  //                          .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  //                          .hps_io_gpio_inst_GPIO61
		output wire [7:0]  led_pio_export,                        //                   led_pio.export
		output wire [14:0] memory_mem_a,                          //                    memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                          .mem_ba
		output wire        memory_mem_ck,                         //                          .mem_ck
		output wire        memory_mem_ck_n,                       //                          .mem_ck_n
		output wire        memory_mem_cke,                        //                          .mem_cke
		output wire        memory_mem_cs_n,                       //                          .mem_cs_n
		output wire        memory_mem_ras_n,                      //                          .mem_ras_n
		output wire        memory_mem_cas_n,                      //                          .mem_cas_n
		output wire        memory_mem_we_n,                       //                          .mem_we_n
		output wire        memory_mem_reset_n,                    //                          .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //                          .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //                          .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //                          .mem_dqs_n
		output wire        memory_mem_odt,                        //                          .mem_odt
		output wire [3:0]  memory_mem_dm,                         //                          .mem_dm
		input  wire        memory_oct_rzqin,                      //                          .oct_rzqin
		input  wire        reset_reset_n                          //                     reset.reset_n
	);

	wire    [1:0] axi_bridge_for_acp_128_0_m0_awburst;                           // axi_bridge_for_acp_128_0:axm_m0_awburst -> hps_0:f2h_AWBURST
	wire    [3:0] axi_bridge_for_acp_128_0_m0_arlen;                             // axi_bridge_for_acp_128_0:axm_m0_arlen -> hps_0:f2h_ARLEN
	wire    [4:0] axi_bridge_for_acp_128_0_m0_awuser;                            // axi_bridge_for_acp_128_0:axm_m0_awuser -> hps_0:f2h_AWUSER
	wire          axi_bridge_for_acp_128_0_m0_wready;                            // hps_0:f2h_WREADY -> axi_bridge_for_acp_128_0:axm_m0_wready
	wire   [15:0] axi_bridge_for_acp_128_0_m0_wstrb;                             // axi_bridge_for_acp_128_0:axm_m0_wstrb -> hps_0:f2h_WSTRB
	wire    [7:0] axi_bridge_for_acp_128_0_m0_rid;                               // hps_0:f2h_RID -> axi_bridge_for_acp_128_0:axm_m0_rid
	wire          axi_bridge_for_acp_128_0_m0_rready;                            // axi_bridge_for_acp_128_0:axm_m0_rready -> hps_0:f2h_RREADY
	wire    [3:0] axi_bridge_for_acp_128_0_m0_awlen;                             // axi_bridge_for_acp_128_0:axm_m0_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] axi_bridge_for_acp_128_0_m0_wid;                               // axi_bridge_for_acp_128_0:axm_m0_wid -> hps_0:f2h_WID
	wire    [3:0] axi_bridge_for_acp_128_0_m0_arcache;                           // axi_bridge_for_acp_128_0:axm_m0_arcache -> hps_0:f2h_ARCACHE
	wire   [31:0] axi_bridge_for_acp_128_0_m0_araddr;                            // axi_bridge_for_acp_128_0:axm_m0_araddr -> hps_0:f2h_ARADDR
	wire          axi_bridge_for_acp_128_0_m0_wvalid;                            // axi_bridge_for_acp_128_0:axm_m0_wvalid -> hps_0:f2h_WVALID
	wire    [2:0] axi_bridge_for_acp_128_0_m0_arprot;                            // axi_bridge_for_acp_128_0:axm_m0_arprot -> hps_0:f2h_ARPROT
	wire          axi_bridge_for_acp_128_0_m0_arvalid;                           // axi_bridge_for_acp_128_0:axm_m0_arvalid -> hps_0:f2h_ARVALID
	wire    [2:0] axi_bridge_for_acp_128_0_m0_awprot;                            // axi_bridge_for_acp_128_0:axm_m0_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] axi_bridge_for_acp_128_0_m0_wdata;                             // axi_bridge_for_acp_128_0:axm_m0_wdata -> hps_0:f2h_WDATA
	wire    [7:0] axi_bridge_for_acp_128_0_m0_arid;                              // axi_bridge_for_acp_128_0:axm_m0_arid -> hps_0:f2h_ARID
	wire    [3:0] axi_bridge_for_acp_128_0_m0_awcache;                           // axi_bridge_for_acp_128_0:axm_m0_awcache -> hps_0:f2h_AWCACHE
	wire    [1:0] axi_bridge_for_acp_128_0_m0_arlock;                            // axi_bridge_for_acp_128_0:axm_m0_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] axi_bridge_for_acp_128_0_m0_awlock;                            // axi_bridge_for_acp_128_0:axm_m0_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] axi_bridge_for_acp_128_0_m0_awaddr;                            // axi_bridge_for_acp_128_0:axm_m0_awaddr -> hps_0:f2h_AWADDR
	wire          axi_bridge_for_acp_128_0_m0_arready;                           // hps_0:f2h_ARREADY -> axi_bridge_for_acp_128_0:axm_m0_arready
	wire    [1:0] axi_bridge_for_acp_128_0_m0_bresp;                             // hps_0:f2h_BRESP -> axi_bridge_for_acp_128_0:axm_m0_bresp
	wire  [127:0] axi_bridge_for_acp_128_0_m0_rdata;                             // hps_0:f2h_RDATA -> axi_bridge_for_acp_128_0:axm_m0_rdata
	wire    [1:0] axi_bridge_for_acp_128_0_m0_arburst;                           // axi_bridge_for_acp_128_0:axm_m0_arburst -> hps_0:f2h_ARBURST
	wire          axi_bridge_for_acp_128_0_m0_awready;                           // hps_0:f2h_AWREADY -> axi_bridge_for_acp_128_0:axm_m0_awready
	wire    [2:0] axi_bridge_for_acp_128_0_m0_arsize;                            // axi_bridge_for_acp_128_0:axm_m0_arsize -> hps_0:f2h_ARSIZE
	wire          axi_bridge_for_acp_128_0_m0_bready;                            // axi_bridge_for_acp_128_0:axm_m0_bready -> hps_0:f2h_BREADY
	wire          axi_bridge_for_acp_128_0_m0_rlast;                             // hps_0:f2h_RLAST -> axi_bridge_for_acp_128_0:axm_m0_rlast
	wire          axi_bridge_for_acp_128_0_m0_wlast;                             // axi_bridge_for_acp_128_0:axm_m0_wlast -> hps_0:f2h_WLAST
	wire    [1:0] axi_bridge_for_acp_128_0_m0_rresp;                             // hps_0:f2h_RRESP -> axi_bridge_for_acp_128_0:axm_m0_rresp
	wire    [7:0] axi_bridge_for_acp_128_0_m0_awid;                              // axi_bridge_for_acp_128_0:axm_m0_awid -> hps_0:f2h_AWID
	wire    [7:0] axi_bridge_for_acp_128_0_m0_bid;                               // hps_0:f2h_BID -> axi_bridge_for_acp_128_0:axm_m0_bid
	wire          axi_bridge_for_acp_128_0_m0_bvalid;                            // hps_0:f2h_BVALID -> axi_bridge_for_acp_128_0:axm_m0_bvalid
	wire    [4:0] axi_bridge_for_acp_128_0_m0_aruser;                            // axi_bridge_for_acp_128_0:axm_m0_aruser -> hps_0:f2h_ARUSER
	wire    [2:0] axi_bridge_for_acp_128_0_m0_awsize;                            // axi_bridge_for_acp_128_0:axm_m0_awsize -> hps_0:f2h_AWSIZE
	wire          axi_bridge_for_acp_128_0_m0_awvalid;                           // axi_bridge_for_acp_128_0:axm_m0_awvalid -> hps_0:f2h_AWVALID
	wire          axi_bridge_for_acp_128_0_m0_rvalid;                            // hps_0:f2h_RVALID -> axi_bridge_for_acp_128_0:axm_m0_rvalid
	wire          hps_0_h2f_user0_clock_clk;                                     // hps_0:h2f_user0_clk -> [axi_bridge_for_acp_128_0:clk, fft_ddr_bridge:clk, fft_sub:clk_clk, hps_0:f2h_axi_clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, mm_interconnect_0:hps_0_h2f_user0_clock_clk, mm_interconnect_3:hps_0_h2f_user0_clock_clk, mm_interconnect_6:hps_0_h2f_user0_clock_clk, rst_controller:clk]
	wire          fft_ddr_bridge_expanded_master_waitrequest;                    // mm_interconnect_0:fft_ddr_bridge_expanded_master_waitrequest -> fft_ddr_bridge:avm_m0_waitrequest
	wire  [127:0] fft_ddr_bridge_expanded_master_readdata;                       // mm_interconnect_0:fft_ddr_bridge_expanded_master_readdata -> fft_ddr_bridge:avm_m0_readdata
	wire   [31:0] fft_ddr_bridge_expanded_master_address;                        // fft_ddr_bridge:avm_m0_address -> mm_interconnect_0:fft_ddr_bridge_expanded_master_address
	wire          fft_ddr_bridge_expanded_master_read;                           // fft_ddr_bridge:avm_m0_read -> mm_interconnect_0:fft_ddr_bridge_expanded_master_read
	wire   [15:0] fft_ddr_bridge_expanded_master_byteenable;                     // fft_ddr_bridge:avm_m0_byteenable -> mm_interconnect_0:fft_ddr_bridge_expanded_master_byteenable
	wire          fft_ddr_bridge_expanded_master_readdatavalid;                  // mm_interconnect_0:fft_ddr_bridge_expanded_master_readdatavalid -> fft_ddr_bridge:avm_m0_readdatavalid
	wire          fft_ddr_bridge_expanded_master_write;                          // fft_ddr_bridge:avm_m0_write -> mm_interconnect_0:fft_ddr_bridge_expanded_master_write
	wire  [127:0] fft_ddr_bridge_expanded_master_writedata;                      // fft_ddr_bridge:avm_m0_writedata -> mm_interconnect_0:fft_ddr_bridge_expanded_master_writedata
	wire    [4:0] fft_ddr_bridge_expanded_master_burstcount;                     // fft_ddr_bridge:avm_m0_burstcount -> mm_interconnect_0:fft_ddr_bridge_expanded_master_burstcount
	wire    [1:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awburst;         // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awburst -> axi_bridge_for_acp_128_0:axs_s0_awburst
	wire    [4:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awuser;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awuser -> axi_bridge_for_acp_128_0:axs_s0_awuser
	wire    [3:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlen;           // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arlen -> axi_bridge_for_acp_128_0:axs_s0_arlen
	wire   [15:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wstrb;           // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wstrb -> axi_bridge_for_acp_128_0:axs_s0_wstrb
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wready;          // axi_bridge_for_acp_128_0:axs_s0_wready -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wready
	wire    [7:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rid;             // axi_bridge_for_acp_128_0:axs_s0_rid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rid
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rready;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rready -> axi_bridge_for_acp_128_0:axs_s0_rready
	wire    [3:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlen;           // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awlen -> axi_bridge_for_acp_128_0:axs_s0_awlen
	wire    [7:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wid;             // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wid -> axi_bridge_for_acp_128_0:axs_s0_wid
	wire    [3:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arcache;         // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arcache -> axi_bridge_for_acp_128_0:axs_s0_arcache
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wvalid;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wvalid -> axi_bridge_for_acp_128_0:axs_s0_wvalid
	wire   [31:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_araddr;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_araddr -> axi_bridge_for_acp_128_0:axs_s0_araddr
	wire    [2:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arprot;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arprot -> axi_bridge_for_acp_128_0:axs_s0_arprot
	wire    [2:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awprot;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awprot -> axi_bridge_for_acp_128_0:axs_s0_awprot
	wire  [127:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wdata;           // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wdata -> axi_bridge_for_acp_128_0:axs_s0_wdata
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arvalid;         // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arvalid -> axi_bridge_for_acp_128_0:axs_s0_arvalid
	wire    [3:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awcache;         // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awcache -> axi_bridge_for_acp_128_0:axs_s0_awcache
	wire    [7:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arid;            // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arid -> axi_bridge_for_acp_128_0:axs_s0_arid
	wire    [1:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlock;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arlock -> axi_bridge_for_acp_128_0:axs_s0_arlock
	wire    [1:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlock;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awlock -> axi_bridge_for_acp_128_0:axs_s0_awlock
	wire   [31:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awaddr;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awaddr -> axi_bridge_for_acp_128_0:axs_s0_awaddr
	wire    [1:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bresp;           // axi_bridge_for_acp_128_0:axs_s0_bresp -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bresp
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arready;         // axi_bridge_for_acp_128_0:axs_s0_arready -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arready
	wire  [127:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rdata;           // axi_bridge_for_acp_128_0:axs_s0_rdata -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rdata
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awready;         // axi_bridge_for_acp_128_0:axs_s0_awready -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awready
	wire    [1:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arburst;         // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arburst -> axi_bridge_for_acp_128_0:axs_s0_arburst
	wire    [2:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arsize;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_arsize -> axi_bridge_for_acp_128_0:axs_s0_arsize
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bready;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bready -> axi_bridge_for_acp_128_0:axs_s0_bready
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rlast;           // axi_bridge_for_acp_128_0:axs_s0_rlast -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rlast
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wlast;           // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_wlast -> axi_bridge_for_acp_128_0:axs_s0_wlast
	wire    [1:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rresp;           // axi_bridge_for_acp_128_0:axs_s0_rresp -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rresp
	wire    [7:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awid;            // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awid -> axi_bridge_for_acp_128_0:axs_s0_awid
	wire    [7:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bid;             // axi_bridge_for_acp_128_0:axs_s0_bid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bid
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bvalid;          // axi_bridge_for_acp_128_0:axs_s0_bvalid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_bvalid
	wire    [2:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awsize;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awsize -> axi_bridge_for_acp_128_0:axs_s0_awsize
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awvalid;         // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_awvalid -> axi_bridge_for_acp_128_0:axs_s0_awvalid
	wire    [4:0] mm_interconnect_0_axi_bridge_for_acp_128_0_s0_aruser;          // mm_interconnect_0:axi_bridge_for_acp_128_0_s0_aruser -> axi_bridge_for_acp_128_0:axs_s0_aruser
	wire          mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rvalid;          // axi_bridge_for_acp_128_0:axs_s0_rvalid -> mm_interconnect_0:axi_bridge_for_acp_128_0_s0_rvalid
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                  // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                    // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                    // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                   // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                      // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                   // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                    // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                      // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                  // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                   // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                   // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                   // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                   // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                    // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                  // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                  // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                     // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                   // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                   // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                   // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                    // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                  // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                  // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                  // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                   // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                   // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                    // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                     // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                      // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                   // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                   // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                  // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                   // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          mm_interconnect_1_onchip_memory2_0_s1_chipselect;              // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;                // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire   [12:0] mm_interconnect_1_onchip_memory2_0_s1_address;                 // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire    [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;              // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_1_onchip_memory2_0_s1_write;                   // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;               // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_1_onchip_memory2_0_s1_clken;                   // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                               // hps_0:h2f_lw_AWBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                 // hps_0:h2f_lw_ARLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                 // hps_0:h2f_lw_WSTRB -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                // mm_interconnect_2:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                   // mm_interconnect_2:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                // hps_0:h2f_lw_RREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                 // hps_0:h2f_lw_AWLEN -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                   // hps_0:h2f_lw_WID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                               // hps_0:h2f_lw_ARCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                // hps_0:h2f_lw_WVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                // hps_0:h2f_lw_ARADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                // hps_0:h2f_lw_ARPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                // hps_0:h2f_lw_AWPROT -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                 // hps_0:h2f_lw_WDATA -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                               // hps_0:h2f_lw_ARVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                               // hps_0:h2f_lw_AWCACHE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                  // hps_0:h2f_lw_ARID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                // hps_0:h2f_lw_ARLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                // hps_0:h2f_lw_AWLOCK -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                // hps_0:h2f_lw_AWADDR -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                               // mm_interconnect_2:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                               // mm_interconnect_2:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                               // hps_0:h2f_lw_ARBURST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                // hps_0:h2f_lw_ARSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                // hps_0:h2f_lw_BREADY -> mm_interconnect_2:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                 // hps_0:h2f_lw_WLAST -> mm_interconnect_2:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                 // mm_interconnect_2:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                  // hps_0:h2f_lw_AWID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                   // mm_interconnect_2:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                // mm_interconnect_2:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                // hps_0:h2f_lw_AWSIZE -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                               // hps_0:h2f_lw_AWVALID -> mm_interconnect_2:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                // mm_interconnect_2:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] fpga_only_master_master_readdata;                              // mm_interconnect_2:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire          fpga_only_master_master_waitrequest;                           // mm_interconnect_2:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire   [31:0] fpga_only_master_master_address;                               // fpga_only_master:master_address -> mm_interconnect_2:fpga_only_master_master_address
	wire          fpga_only_master_master_read;                                  // fpga_only_master:master_read -> mm_interconnect_2:fpga_only_master_master_read
	wire    [3:0] fpga_only_master_master_byteenable;                            // fpga_only_master:master_byteenable -> mm_interconnect_2:fpga_only_master_master_byteenable
	wire          fpga_only_master_master_readdatavalid;                         // mm_interconnect_2:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire          fpga_only_master_master_write;                                 // fpga_only_master:master_write -> mm_interconnect_2:fpga_only_master_master_write
	wire   [31:0] fpga_only_master_master_writedata;                             // fpga_only_master:master_writedata -> mm_interconnect_2:fpga_only_master_master_writedata
	wire   [31:0] mm_interconnect_2_lw_mm_bridge_s0_readdata;                    // lw_mm_bridge:s0_readdata -> mm_interconnect_2:lw_mm_bridge_s0_readdata
	wire          mm_interconnect_2_lw_mm_bridge_s0_waitrequest;                 // lw_mm_bridge:s0_waitrequest -> mm_interconnect_2:lw_mm_bridge_s0_waitrequest
	wire          mm_interconnect_2_lw_mm_bridge_s0_debugaccess;                 // mm_interconnect_2:lw_mm_bridge_s0_debugaccess -> lw_mm_bridge:s0_debugaccess
	wire   [19:0] mm_interconnect_2_lw_mm_bridge_s0_address;                     // mm_interconnect_2:lw_mm_bridge_s0_address -> lw_mm_bridge:s0_address
	wire          mm_interconnect_2_lw_mm_bridge_s0_read;                        // mm_interconnect_2:lw_mm_bridge_s0_read -> lw_mm_bridge:s0_read
	wire    [3:0] mm_interconnect_2_lw_mm_bridge_s0_byteenable;                  // mm_interconnect_2:lw_mm_bridge_s0_byteenable -> lw_mm_bridge:s0_byteenable
	wire          mm_interconnect_2_lw_mm_bridge_s0_readdatavalid;               // lw_mm_bridge:s0_readdatavalid -> mm_interconnect_2:lw_mm_bridge_s0_readdatavalid
	wire          mm_interconnect_2_lw_mm_bridge_s0_write;                       // mm_interconnect_2:lw_mm_bridge_s0_write -> lw_mm_bridge:s0_write
	wire   [31:0] mm_interconnect_2_lw_mm_bridge_s0_writedata;                   // mm_interconnect_2:lw_mm_bridge_s0_writedata -> lw_mm_bridge:s0_writedata
	wire    [0:0] mm_interconnect_2_lw_mm_bridge_s0_burstcount;                  // mm_interconnect_2:lw_mm_bridge_s0_burstcount -> lw_mm_bridge:s0_burstcount
	wire          lw_mm_bridge_m0_waitrequest;                                   // mm_interconnect_3:lw_mm_bridge_m0_waitrequest -> lw_mm_bridge:m0_waitrequest
	wire   [31:0] lw_mm_bridge_m0_readdata;                                      // mm_interconnect_3:lw_mm_bridge_m0_readdata -> lw_mm_bridge:m0_readdata
	wire          lw_mm_bridge_m0_debugaccess;                                   // lw_mm_bridge:m0_debugaccess -> mm_interconnect_3:lw_mm_bridge_m0_debugaccess
	wire   [19:0] lw_mm_bridge_m0_address;                                       // lw_mm_bridge:m0_address -> mm_interconnect_3:lw_mm_bridge_m0_address
	wire          lw_mm_bridge_m0_read;                                          // lw_mm_bridge:m0_read -> mm_interconnect_3:lw_mm_bridge_m0_read
	wire    [3:0] lw_mm_bridge_m0_byteenable;                                    // lw_mm_bridge:m0_byteenable -> mm_interconnect_3:lw_mm_bridge_m0_byteenable
	wire          lw_mm_bridge_m0_readdatavalid;                                 // mm_interconnect_3:lw_mm_bridge_m0_readdatavalid -> lw_mm_bridge:m0_readdatavalid
	wire   [31:0] lw_mm_bridge_m0_writedata;                                     // lw_mm_bridge:m0_writedata -> mm_interconnect_3:lw_mm_bridge_m0_writedata
	wire          lw_mm_bridge_m0_write;                                         // lw_mm_bridge:m0_write -> mm_interconnect_3:lw_mm_bridge_m0_write
	wire    [0:0] lw_mm_bridge_m0_burstcount;                                    // lw_mm_bridge:m0_burstcount -> mm_interconnect_3:lw_mm_bridge_m0_burstcount
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_3:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_3_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_3:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_3:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_3_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_3:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_3:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_3_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_3:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_3_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_3:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata;     // intr_capturer_0:rddata -> mm_interconnect_3:intr_capturer_0_avalon_slave_0_readdata
	wire    [0:0] mm_interconnect_3_intr_capturer_0_avalon_slave_0_address;      // mm_interconnect_3:intr_capturer_0_avalon_slave_0_address -> intr_capturer_0:addr
	wire          mm_interconnect_3_intr_capturer_0_avalon_slave_0_read;         // mm_interconnect_3:intr_capturer_0_avalon_slave_0_read -> intr_capturer_0:read
	wire   [31:0] mm_interconnect_3_sysid_qsys_control_slave_readdata;           // sysid_qsys:readdata -> mm_interconnect_3:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_3_sysid_qsys_control_slave_address;            // mm_interconnect_3:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [63:0] mm_interconnect_3_chip_id_read_mm_0_s0_readdata;               // chip_id_read_mm_0:avs_s0_readdata -> mm_interconnect_3:chip_id_read_mm_0_s0_readdata
	wire          mm_interconnect_3_chip_id_read_mm_0_s0_read;                   // mm_interconnect_3:chip_id_read_mm_0_s0_read -> chip_id_read_mm_0:avs_s0_read
	wire   [31:0] mm_interconnect_3_fft_sub_s0_readdata;                         // fft_sub:s0_readdata -> mm_interconnect_3:fft_sub_s0_readdata
	wire          mm_interconnect_3_fft_sub_s0_waitrequest;                      // fft_sub:s0_waitrequest -> mm_interconnect_3:fft_sub_s0_waitrequest
	wire          mm_interconnect_3_fft_sub_s0_debugaccess;                      // mm_interconnect_3:fft_sub_s0_debugaccess -> fft_sub:s0_debugaccess
	wire   [18:0] mm_interconnect_3_fft_sub_s0_address;                          // mm_interconnect_3:fft_sub_s0_address -> fft_sub:s0_address
	wire          mm_interconnect_3_fft_sub_s0_read;                             // mm_interconnect_3:fft_sub_s0_read -> fft_sub:s0_read
	wire    [3:0] mm_interconnect_3_fft_sub_s0_byteenable;                       // mm_interconnect_3:fft_sub_s0_byteenable -> fft_sub:s0_byteenable
	wire          mm_interconnect_3_fft_sub_s0_readdatavalid;                    // fft_sub:s0_readdatavalid -> mm_interconnect_3:fft_sub_s0_readdatavalid
	wire          mm_interconnect_3_fft_sub_s0_write;                            // mm_interconnect_3:fft_sub_s0_write -> fft_sub:s0_write
	wire   [31:0] mm_interconnect_3_fft_sub_s0_writedata;                        // mm_interconnect_3:fft_sub_s0_writedata -> fft_sub:s0_writedata
	wire    [0:0] mm_interconnect_3_fft_sub_s0_burstcount;                       // mm_interconnect_3:fft_sub_s0_burstcount -> fft_sub:s0_burstcount
	wire          mm_interconnect_3_led_pio_s1_chipselect;                       // mm_interconnect_3:led_pio_s1_chipselect -> led_pio:chipselect
	wire   [31:0] mm_interconnect_3_led_pio_s1_readdata;                         // led_pio:readdata -> mm_interconnect_3:led_pio_s1_readdata
	wire    [1:0] mm_interconnect_3_led_pio_s1_address;                          // mm_interconnect_3:led_pio_s1_address -> led_pio:address
	wire          mm_interconnect_3_led_pio_s1_write;                            // mm_interconnect_3:led_pio_s1_write -> led_pio:write_n
	wire   [31:0] mm_interconnect_3_led_pio_s1_writedata;                        // mm_interconnect_3:led_pio_s1_writedata -> led_pio:writedata
	wire          mm_interconnect_3_dipsw_pio_s1_chipselect;                     // mm_interconnect_3:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	wire   [31:0] mm_interconnect_3_dipsw_pio_s1_readdata;                       // dipsw_pio:readdata -> mm_interconnect_3:dipsw_pio_s1_readdata
	wire    [1:0] mm_interconnect_3_dipsw_pio_s1_address;                        // mm_interconnect_3:dipsw_pio_s1_address -> dipsw_pio:address
	wire          mm_interconnect_3_dipsw_pio_s1_write;                          // mm_interconnect_3:dipsw_pio_s1_write -> dipsw_pio:write_n
	wire   [31:0] mm_interconnect_3_dipsw_pio_s1_writedata;                      // mm_interconnect_3:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	wire          mm_interconnect_3_button_pio_s1_chipselect;                    // mm_interconnect_3:button_pio_s1_chipselect -> button_pio:chipselect
	wire   [31:0] mm_interconnect_3_button_pio_s1_readdata;                      // button_pio:readdata -> mm_interconnect_3:button_pio_s1_readdata
	wire    [1:0] mm_interconnect_3_button_pio_s1_address;                       // mm_interconnect_3:button_pio_s1_address -> button_pio:address
	wire          mm_interconnect_3_button_pio_s1_write;                         // mm_interconnect_3:button_pio_s1_write -> button_pio:write_n
	wire   [31:0] mm_interconnect_3_button_pio_s1_writedata;                     // mm_interconnect_3:button_pio_s1_writedata -> button_pio:writedata
	wire   [31:0] f2sdram_only_master_master_readdata;                           // mm_interconnect_5:f2sdram_only_master_master_readdata -> f2sdram_only_master:master_readdata
	wire          f2sdram_only_master_master_waitrequest;                        // mm_interconnect_5:f2sdram_only_master_master_waitrequest -> f2sdram_only_master:master_waitrequest
	wire   [31:0] f2sdram_only_master_master_address;                            // f2sdram_only_master:master_address -> mm_interconnect_5:f2sdram_only_master_master_address
	wire          f2sdram_only_master_master_read;                               // f2sdram_only_master:master_read -> mm_interconnect_5:f2sdram_only_master_master_read
	wire    [3:0] f2sdram_only_master_master_byteenable;                         // f2sdram_only_master:master_byteenable -> mm_interconnect_5:f2sdram_only_master_master_byteenable
	wire          f2sdram_only_master_master_readdatavalid;                      // mm_interconnect_5:f2sdram_only_master_master_readdatavalid -> f2sdram_only_master:master_readdatavalid
	wire          f2sdram_only_master_master_write;                              // f2sdram_only_master:master_write -> mm_interconnect_5:f2sdram_only_master_master_write
	wire   [31:0] f2sdram_only_master_master_writedata;                          // f2sdram_only_master:master_writedata -> mm_interconnect_5:f2sdram_only_master_master_writedata
	wire    [1:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awburst;               // mm_interconnect_5:hps_0_f2h_sdram0_data_awburst -> hps_0:f2h_sdram0_AWBURST
	wire    [3:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arlen;                 // mm_interconnect_5:hps_0_f2h_sdram0_data_arlen -> hps_0:f2h_sdram0_ARLEN
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_wstrb;                 // mm_interconnect_5:hps_0_f2h_sdram0_data_wstrb -> hps_0:f2h_sdram0_WSTRB
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_wready;                // hps_0:f2h_sdram0_WREADY -> mm_interconnect_5:hps_0_f2h_sdram0_data_wready
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_rid;                   // hps_0:f2h_sdram0_RID -> mm_interconnect_5:hps_0_f2h_sdram0_data_rid
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_rready;                // mm_interconnect_5:hps_0_f2h_sdram0_data_rready -> hps_0:f2h_sdram0_RREADY
	wire    [3:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awlen;                 // mm_interconnect_5:hps_0_f2h_sdram0_data_awlen -> hps_0:f2h_sdram0_AWLEN
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_wid;                   // mm_interconnect_5:hps_0_f2h_sdram0_data_wid -> hps_0:f2h_sdram0_WID
	wire    [3:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arcache;               // mm_interconnect_5:hps_0_f2h_sdram0_data_arcache -> hps_0:f2h_sdram0_ARCACHE
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_wvalid;                // mm_interconnect_5:hps_0_f2h_sdram0_data_wvalid -> hps_0:f2h_sdram0_WVALID
	wire   [31:0] mm_interconnect_5_hps_0_f2h_sdram0_data_araddr;                // mm_interconnect_5:hps_0_f2h_sdram0_data_araddr -> hps_0:f2h_sdram0_ARADDR
	wire    [2:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arprot;                // mm_interconnect_5:hps_0_f2h_sdram0_data_arprot -> hps_0:f2h_sdram0_ARPROT
	wire    [2:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awprot;                // mm_interconnect_5:hps_0_f2h_sdram0_data_awprot -> hps_0:f2h_sdram0_AWPROT
	wire   [63:0] mm_interconnect_5_hps_0_f2h_sdram0_data_wdata;                 // mm_interconnect_5:hps_0_f2h_sdram0_data_wdata -> hps_0:f2h_sdram0_WDATA
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_arvalid;               // mm_interconnect_5:hps_0_f2h_sdram0_data_arvalid -> hps_0:f2h_sdram0_ARVALID
	wire    [3:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awcache;               // mm_interconnect_5:hps_0_f2h_sdram0_data_awcache -> hps_0:f2h_sdram0_AWCACHE
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arid;                  // mm_interconnect_5:hps_0_f2h_sdram0_data_arid -> hps_0:f2h_sdram0_ARID
	wire    [1:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arlock;                // mm_interconnect_5:hps_0_f2h_sdram0_data_arlock -> hps_0:f2h_sdram0_ARLOCK
	wire    [1:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awlock;                // mm_interconnect_5:hps_0_f2h_sdram0_data_awlock -> hps_0:f2h_sdram0_AWLOCK
	wire   [31:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awaddr;                // mm_interconnect_5:hps_0_f2h_sdram0_data_awaddr -> hps_0:f2h_sdram0_AWADDR
	wire    [1:0] mm_interconnect_5_hps_0_f2h_sdram0_data_bresp;                 // hps_0:f2h_sdram0_BRESP -> mm_interconnect_5:hps_0_f2h_sdram0_data_bresp
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_arready;               // hps_0:f2h_sdram0_ARREADY -> mm_interconnect_5:hps_0_f2h_sdram0_data_arready
	wire   [63:0] mm_interconnect_5_hps_0_f2h_sdram0_data_rdata;                 // hps_0:f2h_sdram0_RDATA -> mm_interconnect_5:hps_0_f2h_sdram0_data_rdata
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_awready;               // hps_0:f2h_sdram0_AWREADY -> mm_interconnect_5:hps_0_f2h_sdram0_data_awready
	wire    [1:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arburst;               // mm_interconnect_5:hps_0_f2h_sdram0_data_arburst -> hps_0:f2h_sdram0_ARBURST
	wire    [2:0] mm_interconnect_5_hps_0_f2h_sdram0_data_arsize;                // mm_interconnect_5:hps_0_f2h_sdram0_data_arsize -> hps_0:f2h_sdram0_ARSIZE
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_bready;                // mm_interconnect_5:hps_0_f2h_sdram0_data_bready -> hps_0:f2h_sdram0_BREADY
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_rlast;                 // hps_0:f2h_sdram0_RLAST -> mm_interconnect_5:hps_0_f2h_sdram0_data_rlast
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_wlast;                 // mm_interconnect_5:hps_0_f2h_sdram0_data_wlast -> hps_0:f2h_sdram0_WLAST
	wire    [1:0] mm_interconnect_5_hps_0_f2h_sdram0_data_rresp;                 // hps_0:f2h_sdram0_RRESP -> mm_interconnect_5:hps_0_f2h_sdram0_data_rresp
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awid;                  // mm_interconnect_5:hps_0_f2h_sdram0_data_awid -> hps_0:f2h_sdram0_AWID
	wire    [7:0] mm_interconnect_5_hps_0_f2h_sdram0_data_bid;                   // hps_0:f2h_sdram0_BID -> mm_interconnect_5:hps_0_f2h_sdram0_data_bid
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_bvalid;                // hps_0:f2h_sdram0_BVALID -> mm_interconnect_5:hps_0_f2h_sdram0_data_bvalid
	wire    [2:0] mm_interconnect_5_hps_0_f2h_sdram0_data_awsize;                // mm_interconnect_5:hps_0_f2h_sdram0_data_awsize -> hps_0:f2h_sdram0_AWSIZE
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_awvalid;               // mm_interconnect_5:hps_0_f2h_sdram0_data_awvalid -> hps_0:f2h_sdram0_AWVALID
	wire          mm_interconnect_5_hps_0_f2h_sdram0_data_rvalid;                // hps_0:f2h_sdram0_RVALID -> mm_interconnect_5:hps_0_f2h_sdram0_data_rvalid
	wire          fft_sub_to_ddr_waitrequest;                                    // mm_interconnect_6:fft_sub_to_ddr_waitrequest -> fft_sub:to_ddr_waitrequest
	wire   [63:0] fft_sub_to_ddr_readdata;                                       // mm_interconnect_6:fft_sub_to_ddr_readdata -> fft_sub:to_ddr_readdata
	wire          fft_sub_to_ddr_debugaccess;                                    // fft_sub:to_ddr_debugaccess -> mm_interconnect_6:fft_sub_to_ddr_debugaccess
	wire   [29:0] fft_sub_to_ddr_address;                                        // fft_sub:to_ddr_address -> mm_interconnect_6:fft_sub_to_ddr_address
	wire          fft_sub_to_ddr_read;                                           // fft_sub:to_ddr_read -> mm_interconnect_6:fft_sub_to_ddr_read
	wire    [7:0] fft_sub_to_ddr_byteenable;                                     // fft_sub:to_ddr_byteenable -> mm_interconnect_6:fft_sub_to_ddr_byteenable
	wire          fft_sub_to_ddr_readdatavalid;                                  // mm_interconnect_6:fft_sub_to_ddr_readdatavalid -> fft_sub:to_ddr_readdatavalid
	wire   [63:0] fft_sub_to_ddr_writedata;                                      // fft_sub:to_ddr_writedata -> mm_interconnect_6:fft_sub_to_ddr_writedata
	wire          fft_sub_to_ddr_write;                                          // fft_sub:to_ddr_write -> mm_interconnect_6:fft_sub_to_ddr_write
	wire    [5:0] fft_sub_to_ddr_burstcount;                                     // fft_sub:to_ddr_burstcount -> mm_interconnect_6:fft_sub_to_ddr_burstcount
	wire  [127:0] mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdata;      // fft_ddr_bridge:avs_s0_readdata -> mm_interconnect_6:fft_ddr_bridge_windowed_slave_readdata
	wire          mm_interconnect_6_fft_ddr_bridge_windowed_slave_waitrequest;   // fft_ddr_bridge:avs_s0_waitrequest -> mm_interconnect_6:fft_ddr_bridge_windowed_slave_waitrequest
	wire   [25:0] mm_interconnect_6_fft_ddr_bridge_windowed_slave_address;       // mm_interconnect_6:fft_ddr_bridge_windowed_slave_address -> fft_ddr_bridge:avs_s0_address
	wire          mm_interconnect_6_fft_ddr_bridge_windowed_slave_read;          // mm_interconnect_6:fft_ddr_bridge_windowed_slave_read -> fft_ddr_bridge:avs_s0_read
	wire   [15:0] mm_interconnect_6_fft_ddr_bridge_windowed_slave_byteenable;    // mm_interconnect_6:fft_ddr_bridge_windowed_slave_byteenable -> fft_ddr_bridge:avs_s0_byteenable
	wire          mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdatavalid; // fft_ddr_bridge:avs_s0_readdatavalid -> mm_interconnect_6:fft_ddr_bridge_windowed_slave_readdatavalid
	wire          mm_interconnect_6_fft_ddr_bridge_windowed_slave_write;         // mm_interconnect_6:fft_ddr_bridge_windowed_slave_write -> fft_ddr_bridge:avs_s0_write
	wire  [127:0] mm_interconnect_6_fft_ddr_bridge_windowed_slave_writedata;     // mm_interconnect_6:fft_ddr_bridge_windowed_slave_writedata -> fft_ddr_bridge:avs_s0_writedata
	wire    [4:0] mm_interconnect_6_fft_ddr_bridge_windowed_slave_burstcount;    // mm_interconnect_6:fft_ddr_bridge_windowed_slave_burstcount -> fft_ddr_bridge:avs_s0_burstcount
	wire   [31:0] hps_0_f2h_irq0_irq;                                            // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                            // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire   [31:0] intr_capturer_0_interrupt_receiver_irq;                        // irq_mapper_002:sender_irq -> intr_capturer_0:interrupt_in
	wire          irq_mapper_002_receiver3_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper_002:receiver3_irq
	wire          irq_mapper_002_receiver4_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper_002:receiver4_irq
	wire          irq_mapper_002_receiver5_irq;                                  // irq_synchronizer_002:sender_irq -> irq_mapper_002:receiver5_irq
	wire          irq_mapper_receiver2_irq;                                      // button_pio:irq -> [irq_mapper:receiver2_irq, irq_mapper_002:receiver2_irq]
	wire          irq_mapper_receiver1_irq;                                      // dipsw_pio:irq -> [irq_mapper:receiver1_irq, irq_mapper_002:receiver1_irq]
	wire          irq_mapper_receiver3_irq;                                      // fft_sub:sgdma_from_fft_csr_irq_irq -> [irq_mapper:receiver3_irq, irq_synchronizer:receiver_irq]
	wire          irq_mapper_receiver4_irq;                                      // fft_sub:sgdma_from_ram_csr_irq_irq -> [irq_mapper:receiver4_irq, irq_synchronizer_001:receiver_irq]
	wire          irq_mapper_receiver5_irq;                                      // fft_sub:sgdma_to_fft_csr_irq_irq -> [irq_mapper:receiver5_irq, irq_synchronizer_002:receiver_irq]
	wire          irq_mapper_receiver0_irq;                                      // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq]
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [axi_bridge_for_acp_128_0:reset, fft_ddr_bridge:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, mm_interconnect_0:fft_ddr_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_3:fft_sub_reset_reset_bridge_in_reset_reset, mm_interconnect_3:fft_sub_s0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_6:fft_ddr_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_6:fft_sub_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [button_pio:reset_n, chip_id_read_mm_0:reset, dipsw_pio:reset_n, intr_capturer_0:rst_n, irq_mapper_002:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart:rst_n, led_pio:reset_n, lw_mm_bridge:reset, mm_interconnect_1:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_2:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:lw_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_3:lw_mm_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_5:f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_5:f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys:reset_n]
	wire          rst_controller_001_reset_out_reset_req;                        // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> [mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_5:hps_0_f2h_sdram0_data_agent_reset_sink_reset_bridge_in_reset_reset]

	axi_bridge_for_acp_128 axi_bridge_for_acp_128_0 (
		.clk            (hps_0_h2f_user0_clock_clk),                             // clock.clk
		.reset          (rst_controller_reset_out_reset),                        // reset.reset
		.axm_m0_araddr  (axi_bridge_for_acp_128_0_m0_araddr),                    //    m0.araddr
		.axm_m0_arburst (axi_bridge_for_acp_128_0_m0_arburst),                   //      .arburst
		.axm_m0_arcache (axi_bridge_for_acp_128_0_m0_arcache),                   //      .arcache
		.axm_m0_arid    (axi_bridge_for_acp_128_0_m0_arid),                      //      .arid
		.axm_m0_arlen   (axi_bridge_for_acp_128_0_m0_arlen),                     //      .arlen
		.axm_m0_arlock  (axi_bridge_for_acp_128_0_m0_arlock),                    //      .arlock
		.axm_m0_arprot  (axi_bridge_for_acp_128_0_m0_arprot),                    //      .arprot
		.axm_m0_arready (axi_bridge_for_acp_128_0_m0_arready),                   //      .arready
		.axm_m0_arsize  (axi_bridge_for_acp_128_0_m0_arsize),                    //      .arsize
		.axm_m0_aruser  (axi_bridge_for_acp_128_0_m0_aruser),                    //      .aruser
		.axm_m0_arvalid (axi_bridge_for_acp_128_0_m0_arvalid),                   //      .arvalid
		.axm_m0_awaddr  (axi_bridge_for_acp_128_0_m0_awaddr),                    //      .awaddr
		.axm_m0_awburst (axi_bridge_for_acp_128_0_m0_awburst),                   //      .awburst
		.axm_m0_awcache (axi_bridge_for_acp_128_0_m0_awcache),                   //      .awcache
		.axm_m0_awid    (axi_bridge_for_acp_128_0_m0_awid),                      //      .awid
		.axm_m0_awlen   (axi_bridge_for_acp_128_0_m0_awlen),                     //      .awlen
		.axm_m0_awlock  (axi_bridge_for_acp_128_0_m0_awlock),                    //      .awlock
		.axm_m0_awprot  (axi_bridge_for_acp_128_0_m0_awprot),                    //      .awprot
		.axm_m0_awready (axi_bridge_for_acp_128_0_m0_awready),                   //      .awready
		.axm_m0_awsize  (axi_bridge_for_acp_128_0_m0_awsize),                    //      .awsize
		.axm_m0_awuser  (axi_bridge_for_acp_128_0_m0_awuser),                    //      .awuser
		.axm_m0_awvalid (axi_bridge_for_acp_128_0_m0_awvalid),                   //      .awvalid
		.axm_m0_bid     (axi_bridge_for_acp_128_0_m0_bid),                       //      .bid
		.axm_m0_bready  (axi_bridge_for_acp_128_0_m0_bready),                    //      .bready
		.axm_m0_bresp   (axi_bridge_for_acp_128_0_m0_bresp),                     //      .bresp
		.axm_m0_bvalid  (axi_bridge_for_acp_128_0_m0_bvalid),                    //      .bvalid
		.axm_m0_rdata   (axi_bridge_for_acp_128_0_m0_rdata),                     //      .rdata
		.axm_m0_rid     (axi_bridge_for_acp_128_0_m0_rid),                       //      .rid
		.axm_m0_rlast   (axi_bridge_for_acp_128_0_m0_rlast),                     //      .rlast
		.axm_m0_rready  (axi_bridge_for_acp_128_0_m0_rready),                    //      .rready
		.axm_m0_rresp   (axi_bridge_for_acp_128_0_m0_rresp),                     //      .rresp
		.axm_m0_rvalid  (axi_bridge_for_acp_128_0_m0_rvalid),                    //      .rvalid
		.axm_m0_wdata   (axi_bridge_for_acp_128_0_m0_wdata),                     //      .wdata
		.axm_m0_wid     (axi_bridge_for_acp_128_0_m0_wid),                       //      .wid
		.axm_m0_wlast   (axi_bridge_for_acp_128_0_m0_wlast),                     //      .wlast
		.axm_m0_wready  (axi_bridge_for_acp_128_0_m0_wready),                    //      .wready
		.axm_m0_wstrb   (axi_bridge_for_acp_128_0_m0_wstrb),                     //      .wstrb
		.axm_m0_wvalid  (axi_bridge_for_acp_128_0_m0_wvalid),                    //      .wvalid
		.axs_s0_araddr  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_araddr),  //    s0.araddr
		.axs_s0_arburst (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arburst), //      .arburst
		.axs_s0_arcache (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arcache), //      .arcache
		.axs_s0_arid    (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arid),    //      .arid
		.axs_s0_arlen   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlen),   //      .arlen
		.axs_s0_arlock  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlock),  //      .arlock
		.axs_s0_arprot  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arprot),  //      .arprot
		.axs_s0_arready (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arready), //      .arready
		.axs_s0_arsize  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arsize),  //      .arsize
		.axs_s0_aruser  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_aruser),  //      .aruser
		.axs_s0_arvalid (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arvalid), //      .arvalid
		.axs_s0_awaddr  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awaddr),  //      .awaddr
		.axs_s0_awburst (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awburst), //      .awburst
		.axs_s0_awcache (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awcache), //      .awcache
		.axs_s0_awid    (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awid),    //      .awid
		.axs_s0_awlen   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlen),   //      .awlen
		.axs_s0_awlock  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlock),  //      .awlock
		.axs_s0_awprot  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awprot),  //      .awprot
		.axs_s0_awready (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awready), //      .awready
		.axs_s0_awsize  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awsize),  //      .awsize
		.axs_s0_awuser  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awuser),  //      .awuser
		.axs_s0_awvalid (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awvalid), //      .awvalid
		.axs_s0_bid     (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bid),     //      .bid
		.axs_s0_bready  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bready),  //      .bready
		.axs_s0_bresp   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bresp),   //      .bresp
		.axs_s0_bvalid  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bvalid),  //      .bvalid
		.axs_s0_rdata   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rdata),   //      .rdata
		.axs_s0_rid     (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rid),     //      .rid
		.axs_s0_rlast   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rlast),   //      .rlast
		.axs_s0_rready  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rready),  //      .rready
		.axs_s0_rresp   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rresp),   //      .rresp
		.axs_s0_rvalid  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rvalid),  //      .rvalid
		.axs_s0_wdata   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wdata),   //      .wdata
		.axs_s0_wid     (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wid),     //      .wid
		.axs_s0_wlast   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wlast),   //      .wlast
		.axs_s0_wready  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wready),  //      .wready
		.axs_s0_wstrb   (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wstrb),   //      .wstrb
		.axs_s0_wvalid  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wvalid)   //      .wvalid
	);

	soc_system_button_pio button_pio (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_3_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	chip_id_read_mm chip_id_read_mm_0 (
		.clk             (clk_clk),                                         // clock.clk
		.reset           (rst_controller_001_reset_out_reset),              // reset.reset
		.avs_s0_read     (mm_interconnect_3_chip_id_read_mm_0_s0_read),     //    s0.read
		.avs_s0_readdata (mm_interconnect_3_chip_id_read_mm_0_s0_readdata), //      .readdata
		.asi_in0_data    (),                                                //   in0.data
		.asi_in0_ready   ()                                                 //      .ready
	);

	soc_system_dipsw_pio dipsw_pio (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_3_dipsw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_dipsw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_dipsw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_dipsw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_dipsw_pio_s1_readdata),   //                    .readdata
		.in_port    (dipsw_pio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) f2sdram_only_master (
		.clk_clk              (clk_clk),                                  //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                           //    clk_reset.reset
		.master_address       (f2sdram_only_master_master_address),       //       master.address
		.master_readdata      (f2sdram_only_master_master_readdata),      //             .readdata
		.master_read          (f2sdram_only_master_master_read),          //             .read
		.master_write         (f2sdram_only_master_master_write),         //             .write
		.master_writedata     (f2sdram_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (f2sdram_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (f2sdram_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (f2sdram_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	altera_address_span_extender #(
		.DATA_WIDTH           (128),
		.BYTEENABLE_WIDTH     (16),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (26),
		.SLAVE_ADDRESS_SHIFT  (4),
		.BURSTCOUNT_WIDTH     (5),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000010000000000000000000000000000000)
	) fft_ddr_bridge (
		.clk                  (hps_0_h2f_user0_clock_clk),                                     //           clock.clk
		.reset                (rst_controller_reset_out_reset),                                //           reset.reset
		.avs_s0_address       (mm_interconnect_6_fft_ddr_bridge_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_6_fft_ddr_bridge_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_6_fft_ddr_bridge_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_6_fft_ddr_bridge_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_6_fft_ddr_bridge_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_6_fft_ddr_bridge_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_6_fft_ddr_bridge_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (fft_ddr_bridge_expanded_master_address),                        // expanded_master.address
		.avm_m0_read          (fft_ddr_bridge_expanded_master_read),                           //                .read
		.avm_m0_waitrequest   (fft_ddr_bridge_expanded_master_waitrequest),                    //                .waitrequest
		.avm_m0_readdata      (fft_ddr_bridge_expanded_master_readdata),                       //                .readdata
		.avm_m0_write         (fft_ddr_bridge_expanded_master_write),                          //                .write
		.avm_m0_writedata     (fft_ddr_bridge_expanded_master_writedata),                      //                .writedata
		.avm_m0_readdatavalid (fft_ddr_bridge_expanded_master_readdatavalid),                  //                .readdatavalid
		.avm_m0_byteenable    (fft_ddr_bridge_expanded_master_byteenable),                     //                .byteenable
		.avm_m0_burstcount    (fft_ddr_bridge_expanded_master_burstcount),                     //                .burstcount
		.avs_cntl_read        (),                                                              //            cntl.read
		.avs_cntl_readdata    (),                                                              //                .readdata
		.avs_cntl_write       (),                                                              //                .write
		.avs_cntl_writedata   (),                                                              //                .writedata
		.avs_cntl_byteenable  (),                                                              //                .byteenable
		.avs_cntl_address     (1'b0)                                                           //     (terminated)
	);

	soc_system_fft_sub fft_sub (
		.clk_clk                    (hps_0_h2f_user0_clock_clk),                  //                    clk.clk
		.reset_reset_n              (reset_reset_n),                              //                  reset.reset_n
		.s0_waitrequest             (mm_interconnect_3_fft_sub_s0_waitrequest),   //                     s0.waitrequest
		.s0_readdata                (mm_interconnect_3_fft_sub_s0_readdata),      //                       .readdata
		.s0_readdatavalid           (mm_interconnect_3_fft_sub_s0_readdatavalid), //                       .readdatavalid
		.s0_burstcount              (mm_interconnect_3_fft_sub_s0_burstcount),    //                       .burstcount
		.s0_writedata               (mm_interconnect_3_fft_sub_s0_writedata),     //                       .writedata
		.s0_address                 (mm_interconnect_3_fft_sub_s0_address),       //                       .address
		.s0_write                   (mm_interconnect_3_fft_sub_s0_write),         //                       .write
		.s0_read                    (mm_interconnect_3_fft_sub_s0_read),          //                       .read
		.s0_byteenable              (mm_interconnect_3_fft_sub_s0_byteenable),    //                       .byteenable
		.s0_debugaccess             (mm_interconnect_3_fft_sub_s0_debugaccess),   //                       .debugaccess
		.sgdma_from_fft_csr_irq_irq (irq_mapper_receiver3_irq),                   // sgdma_from_fft_csr_irq.irq
		.sgdma_from_ram_csr_irq_irq (irq_mapper_receiver4_irq),                   // sgdma_from_ram_csr_irq.irq
		.sgdma_to_fft_csr_irq_irq   (irq_mapper_receiver5_irq),                   //   sgdma_to_fft_csr_irq.irq
		.to_ddr_waitrequest         (fft_sub_to_ddr_waitrequest),                 //                 to_ddr.waitrequest
		.to_ddr_readdata            (fft_sub_to_ddr_readdata),                    //                       .readdata
		.to_ddr_readdatavalid       (fft_sub_to_ddr_readdatavalid),               //                       .readdatavalid
		.to_ddr_burstcount          (fft_sub_to_ddr_burstcount),                  //                       .burstcount
		.to_ddr_writedata           (fft_sub_to_ddr_writedata),                   //                       .writedata
		.to_ddr_address             (fft_sub_to_ddr_address),                     //                       .address
		.to_ddr_write               (fft_sub_to_ddr_write),                       //                       .write
		.to_ddr_read                (fft_sub_to_ddr_read),                        //                       .read
		.to_ddr_byteenable          (fft_sub_to_ddr_byteenable),                  //                       .byteenable
		.to_ddr_debugaccess         (fft_sub_to_ddr_debugaccess)                  //                       .debugaccess
	);

	soc_system_f2sdram_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (clk_clk),                               //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                        //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),                //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),               // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),                //  f2h_warm_reset_req.reset_n
		.h2f_user0_clk            (hps_0_h2f_user0_clock_clk),                       //     h2f_user0_clock.clk
		.h2f_user1_clk            (hps_0_h2f_clk_clk),                               //     h2f_user1_clock.clk
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),            //   f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                                    //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                   //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                   //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                 //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                  //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                 //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                 //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                              //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                   //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                  //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                  //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                   //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),           //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),             //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),             //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),             //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),             //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),             //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),             //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),              //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),           //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),           //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),           //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),             //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),             //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),             //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),               //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),               //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),               //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),               //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),               //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),               //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),              //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),             //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),             //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),              //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),               //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),               //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),               //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),               //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),               //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),               //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),            //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),            //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),            //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),            //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),            //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),            //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                         //           h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                                         //    f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR        (mm_interconnect_5_hps_0_f2h_sdram0_data_araddr),  //     f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN         (mm_interconnect_5_hps_0_f2h_sdram0_data_arlen),   //                    .arlen
		.f2h_sdram0_ARID          (mm_interconnect_5_hps_0_f2h_sdram0_data_arid),    //                    .arid
		.f2h_sdram0_ARSIZE        (mm_interconnect_5_hps_0_f2h_sdram0_data_arsize),  //                    .arsize
		.f2h_sdram0_ARBURST       (mm_interconnect_5_hps_0_f2h_sdram0_data_arburst), //                    .arburst
		.f2h_sdram0_ARLOCK        (mm_interconnect_5_hps_0_f2h_sdram0_data_arlock),  //                    .arlock
		.f2h_sdram0_ARPROT        (mm_interconnect_5_hps_0_f2h_sdram0_data_arprot),  //                    .arprot
		.f2h_sdram0_ARVALID       (mm_interconnect_5_hps_0_f2h_sdram0_data_arvalid), //                    .arvalid
		.f2h_sdram0_ARCACHE       (mm_interconnect_5_hps_0_f2h_sdram0_data_arcache), //                    .arcache
		.f2h_sdram0_AWADDR        (mm_interconnect_5_hps_0_f2h_sdram0_data_awaddr),  //                    .awaddr
		.f2h_sdram0_AWLEN         (mm_interconnect_5_hps_0_f2h_sdram0_data_awlen),   //                    .awlen
		.f2h_sdram0_AWID          (mm_interconnect_5_hps_0_f2h_sdram0_data_awid),    //                    .awid
		.f2h_sdram0_AWSIZE        (mm_interconnect_5_hps_0_f2h_sdram0_data_awsize),  //                    .awsize
		.f2h_sdram0_AWBURST       (mm_interconnect_5_hps_0_f2h_sdram0_data_awburst), //                    .awburst
		.f2h_sdram0_AWLOCK        (mm_interconnect_5_hps_0_f2h_sdram0_data_awlock),  //                    .awlock
		.f2h_sdram0_AWPROT        (mm_interconnect_5_hps_0_f2h_sdram0_data_awprot),  //                    .awprot
		.f2h_sdram0_AWVALID       (mm_interconnect_5_hps_0_f2h_sdram0_data_awvalid), //                    .awvalid
		.f2h_sdram0_AWCACHE       (mm_interconnect_5_hps_0_f2h_sdram0_data_awcache), //                    .awcache
		.f2h_sdram0_BRESP         (mm_interconnect_5_hps_0_f2h_sdram0_data_bresp),   //                    .bresp
		.f2h_sdram0_BID           (mm_interconnect_5_hps_0_f2h_sdram0_data_bid),     //                    .bid
		.f2h_sdram0_BVALID        (mm_interconnect_5_hps_0_f2h_sdram0_data_bvalid),  //                    .bvalid
		.f2h_sdram0_BREADY        (mm_interconnect_5_hps_0_f2h_sdram0_data_bready),  //                    .bready
		.f2h_sdram0_ARREADY       (mm_interconnect_5_hps_0_f2h_sdram0_data_arready), //                    .arready
		.f2h_sdram0_AWREADY       (mm_interconnect_5_hps_0_f2h_sdram0_data_awready), //                    .awready
		.f2h_sdram0_RREADY        (mm_interconnect_5_hps_0_f2h_sdram0_data_rready),  //                    .rready
		.f2h_sdram0_RDATA         (mm_interconnect_5_hps_0_f2h_sdram0_data_rdata),   //                    .rdata
		.f2h_sdram0_RRESP         (mm_interconnect_5_hps_0_f2h_sdram0_data_rresp),   //                    .rresp
		.f2h_sdram0_RLAST         (mm_interconnect_5_hps_0_f2h_sdram0_data_rlast),   //                    .rlast
		.f2h_sdram0_RID           (mm_interconnect_5_hps_0_f2h_sdram0_data_rid),     //                    .rid
		.f2h_sdram0_RVALID        (mm_interconnect_5_hps_0_f2h_sdram0_data_rvalid),  //                    .rvalid
		.f2h_sdram0_WLAST         (mm_interconnect_5_hps_0_f2h_sdram0_data_wlast),   //                    .wlast
		.f2h_sdram0_WVALID        (mm_interconnect_5_hps_0_f2h_sdram0_data_wvalid),  //                    .wvalid
		.f2h_sdram0_WDATA         (mm_interconnect_5_hps_0_f2h_sdram0_data_wdata),   //                    .wdata
		.f2h_sdram0_WSTRB         (mm_interconnect_5_hps_0_f2h_sdram0_data_wstrb),   //                    .wstrb
		.f2h_sdram0_WREADY        (mm_interconnect_5_hps_0_f2h_sdram0_data_wready),  //                    .wready
		.f2h_sdram0_WID           (mm_interconnect_5_hps_0_f2h_sdram0_data_wid),     //                    .wid
		.h2f_axi_clk              (clk_clk),                                         //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                       //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                     //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                      //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                     //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                    //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                     //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                    //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                     //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                    //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                    //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                        //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                      //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                      //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                      //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                     //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                     //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                        //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                      //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                     //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                     //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                       //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                     //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                      //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                     //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                    //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                     //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                    //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                     //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                    //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                    //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                        //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                      //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                      //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                      //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                     //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                     //                    .rready
		.f2h_axi_clk              (hps_0_h2f_user0_clock_clk),                       //       f2h_axi_clock.clk
		.f2h_AWID                 (axi_bridge_for_acp_128_0_m0_awid),                //       f2h_axi_slave.awid
		.f2h_AWADDR               (axi_bridge_for_acp_128_0_m0_awaddr),              //                    .awaddr
		.f2h_AWLEN                (axi_bridge_for_acp_128_0_m0_awlen),               //                    .awlen
		.f2h_AWSIZE               (axi_bridge_for_acp_128_0_m0_awsize),              //                    .awsize
		.f2h_AWBURST              (axi_bridge_for_acp_128_0_m0_awburst),             //                    .awburst
		.f2h_AWLOCK               (axi_bridge_for_acp_128_0_m0_awlock),              //                    .awlock
		.f2h_AWCACHE              (axi_bridge_for_acp_128_0_m0_awcache),             //                    .awcache
		.f2h_AWPROT               (axi_bridge_for_acp_128_0_m0_awprot),              //                    .awprot
		.f2h_AWVALID              (axi_bridge_for_acp_128_0_m0_awvalid),             //                    .awvalid
		.f2h_AWREADY              (axi_bridge_for_acp_128_0_m0_awready),             //                    .awready
		.f2h_AWUSER               (axi_bridge_for_acp_128_0_m0_awuser),              //                    .awuser
		.f2h_WID                  (axi_bridge_for_acp_128_0_m0_wid),                 //                    .wid
		.f2h_WDATA                (axi_bridge_for_acp_128_0_m0_wdata),               //                    .wdata
		.f2h_WSTRB                (axi_bridge_for_acp_128_0_m0_wstrb),               //                    .wstrb
		.f2h_WLAST                (axi_bridge_for_acp_128_0_m0_wlast),               //                    .wlast
		.f2h_WVALID               (axi_bridge_for_acp_128_0_m0_wvalid),              //                    .wvalid
		.f2h_WREADY               (axi_bridge_for_acp_128_0_m0_wready),              //                    .wready
		.f2h_BID                  (axi_bridge_for_acp_128_0_m0_bid),                 //                    .bid
		.f2h_BRESP                (axi_bridge_for_acp_128_0_m0_bresp),               //                    .bresp
		.f2h_BVALID               (axi_bridge_for_acp_128_0_m0_bvalid),              //                    .bvalid
		.f2h_BREADY               (axi_bridge_for_acp_128_0_m0_bready),              //                    .bready
		.f2h_ARID                 (axi_bridge_for_acp_128_0_m0_arid),                //                    .arid
		.f2h_ARADDR               (axi_bridge_for_acp_128_0_m0_araddr),              //                    .araddr
		.f2h_ARLEN                (axi_bridge_for_acp_128_0_m0_arlen),               //                    .arlen
		.f2h_ARSIZE               (axi_bridge_for_acp_128_0_m0_arsize),              //                    .arsize
		.f2h_ARBURST              (axi_bridge_for_acp_128_0_m0_arburst),             //                    .arburst
		.f2h_ARLOCK               (axi_bridge_for_acp_128_0_m0_arlock),              //                    .arlock
		.f2h_ARCACHE              (axi_bridge_for_acp_128_0_m0_arcache),             //                    .arcache
		.f2h_ARPROT               (axi_bridge_for_acp_128_0_m0_arprot),              //                    .arprot
		.f2h_ARVALID              (axi_bridge_for_acp_128_0_m0_arvalid),             //                    .arvalid
		.f2h_ARREADY              (axi_bridge_for_acp_128_0_m0_arready),             //                    .arready
		.f2h_ARUSER               (axi_bridge_for_acp_128_0_m0_aruser),              //                    .aruser
		.f2h_RID                  (axi_bridge_for_acp_128_0_m0_rid),                 //                    .rid
		.f2h_RDATA                (axi_bridge_for_acp_128_0_m0_rdata),               //                    .rdata
		.f2h_RRESP                (axi_bridge_for_acp_128_0_m0_rresp),               //                    .rresp
		.f2h_RLAST                (axi_bridge_for_acp_128_0_m0_rlast),               //                    .rlast
		.f2h_RVALID               (axi_bridge_for_acp_128_0_m0_rvalid),              //                    .rvalid
		.f2h_RREADY               (axi_bridge_for_acp_128_0_m0_rready),              //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                                         //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                    //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                  //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                   //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                  //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                 //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                  //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                 //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                  //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                 //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                 //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                     //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                   //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                   //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                   //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                  //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                  //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                     //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                   //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                  //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                  //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                    //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                  //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                   //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                  //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                 //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                  //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                 //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                  //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                 //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                 //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                     //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                   //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                   //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                   //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                  //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                  //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                              //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                               //            f2h_irq1.irq
	);

	intr_capturer #(
		.NUM_INTR (32)
	) intr_capturer_0 (
		.clk          (clk_clk),                                                   //              clock.clk
		.rst_n        (~rst_controller_001_reset_out_reset),                       //         reset_sink.reset_n
		.addr         (mm_interconnect_3_intr_capturer_0_avalon_slave_0_address),  //     avalon_slave_0.address
		.read         (mm_interconnect_3_intr_capturer_0_avalon_slave_0_read),     //                   .read
		.rddata       (mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata), //                   .readdata
		.interrupt_in (intr_capturer_0_interrupt_receiver_irq)                     // interrupt_receiver.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_3_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_3_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_3_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_3_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_3_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_3_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_3_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	soc_system_led_pio led_pio (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_3_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (20),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) lw_mm_bridge (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),              // reset.reset
		.s0_waitrequest   (mm_interconnect_2_lw_mm_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_2_lw_mm_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_2_lw_mm_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_2_lw_mm_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_2_lw_mm_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_2_lw_mm_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_2_lw_mm_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_2_lw_mm_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_2_lw_mm_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_2_lw_mm_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (lw_mm_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (lw_mm_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (lw_mm_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (lw_mm_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (lw_mm_bridge_m0_writedata),                       //      .writedata
		.m0_address       (lw_mm_bridge_m0_address),                         //      .address
		.m0_write         (lw_mm_bridge_m0_write),                           //      .write
		.m0_read          (lw_mm_bridge_m0_read),                            //      .read
		.m0_byteenable    (lw_mm_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (lw_mm_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                // (terminated)
		.m0_response      (2'b00)                                            // (terminated)
	);

	soc_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_3_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_3_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.axi_bridge_for_acp_128_0_s0_awid                 (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awid),    //                axi_bridge_for_acp_128_0_s0.awid
		.axi_bridge_for_acp_128_0_s0_awaddr               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awaddr),  //                                           .awaddr
		.axi_bridge_for_acp_128_0_s0_awlen                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlen),   //                                           .awlen
		.axi_bridge_for_acp_128_0_s0_awsize               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awsize),  //                                           .awsize
		.axi_bridge_for_acp_128_0_s0_awburst              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awburst), //                                           .awburst
		.axi_bridge_for_acp_128_0_s0_awlock               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awlock),  //                                           .awlock
		.axi_bridge_for_acp_128_0_s0_awcache              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awcache), //                                           .awcache
		.axi_bridge_for_acp_128_0_s0_awprot               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awprot),  //                                           .awprot
		.axi_bridge_for_acp_128_0_s0_awuser               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awuser),  //                                           .awuser
		.axi_bridge_for_acp_128_0_s0_awvalid              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awvalid), //                                           .awvalid
		.axi_bridge_for_acp_128_0_s0_awready              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_awready), //                                           .awready
		.axi_bridge_for_acp_128_0_s0_wid                  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wid),     //                                           .wid
		.axi_bridge_for_acp_128_0_s0_wdata                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wdata),   //                                           .wdata
		.axi_bridge_for_acp_128_0_s0_wstrb                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wstrb),   //                                           .wstrb
		.axi_bridge_for_acp_128_0_s0_wlast                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wlast),   //                                           .wlast
		.axi_bridge_for_acp_128_0_s0_wvalid               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wvalid),  //                                           .wvalid
		.axi_bridge_for_acp_128_0_s0_wready               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_wready),  //                                           .wready
		.axi_bridge_for_acp_128_0_s0_bid                  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bid),     //                                           .bid
		.axi_bridge_for_acp_128_0_s0_bresp                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bresp),   //                                           .bresp
		.axi_bridge_for_acp_128_0_s0_bvalid               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bvalid),  //                                           .bvalid
		.axi_bridge_for_acp_128_0_s0_bready               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_bready),  //                                           .bready
		.axi_bridge_for_acp_128_0_s0_arid                 (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arid),    //                                           .arid
		.axi_bridge_for_acp_128_0_s0_araddr               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_araddr),  //                                           .araddr
		.axi_bridge_for_acp_128_0_s0_arlen                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlen),   //                                           .arlen
		.axi_bridge_for_acp_128_0_s0_arsize               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arsize),  //                                           .arsize
		.axi_bridge_for_acp_128_0_s0_arburst              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arburst), //                                           .arburst
		.axi_bridge_for_acp_128_0_s0_arlock               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arlock),  //                                           .arlock
		.axi_bridge_for_acp_128_0_s0_arcache              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arcache), //                                           .arcache
		.axi_bridge_for_acp_128_0_s0_arprot               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arprot),  //                                           .arprot
		.axi_bridge_for_acp_128_0_s0_aruser               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_aruser),  //                                           .aruser
		.axi_bridge_for_acp_128_0_s0_arvalid              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arvalid), //                                           .arvalid
		.axi_bridge_for_acp_128_0_s0_arready              (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_arready), //                                           .arready
		.axi_bridge_for_acp_128_0_s0_rid                  (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rid),     //                                           .rid
		.axi_bridge_for_acp_128_0_s0_rdata                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rdata),   //                                           .rdata
		.axi_bridge_for_acp_128_0_s0_rresp                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rresp),   //                                           .rresp
		.axi_bridge_for_acp_128_0_s0_rlast                (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rlast),   //                                           .rlast
		.axi_bridge_for_acp_128_0_s0_rvalid               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rvalid),  //                                           .rvalid
		.axi_bridge_for_acp_128_0_s0_rready               (mm_interconnect_0_axi_bridge_for_acp_128_0_s0_rready),  //                                           .rready
		.hps_0_h2f_user0_clock_clk                        (hps_0_h2f_user0_clock_clk),                             //                      hps_0_h2f_user0_clock.clk
		.fft_ddr_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // fft_ddr_bridge_reset_reset_bridge_in_reset.reset
		.fft_ddr_bridge_expanded_master_address           (fft_ddr_bridge_expanded_master_address),                //             fft_ddr_bridge_expanded_master.address
		.fft_ddr_bridge_expanded_master_waitrequest       (fft_ddr_bridge_expanded_master_waitrequest),            //                                           .waitrequest
		.fft_ddr_bridge_expanded_master_burstcount        (fft_ddr_bridge_expanded_master_burstcount),             //                                           .burstcount
		.fft_ddr_bridge_expanded_master_byteenable        (fft_ddr_bridge_expanded_master_byteenable),             //                                           .byteenable
		.fft_ddr_bridge_expanded_master_read              (fft_ddr_bridge_expanded_master_read),                   //                                           .read
		.fft_ddr_bridge_expanded_master_readdata          (fft_ddr_bridge_expanded_master_readdata),               //                                           .readdata
		.fft_ddr_bridge_expanded_master_readdatavalid     (fft_ddr_bridge_expanded_master_readdatavalid),          //                                           .readdatavalid
		.fft_ddr_bridge_expanded_master_write             (fft_ddr_bridge_expanded_master_write),                  //                                           .write
		.fft_ddr_bridge_expanded_master_writedata         (fft_ddr_bridge_expanded_master_writedata)               //                                           .writedata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                        //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                      //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                       //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                      //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                     //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                      //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                     //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                      //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                     //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                     //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                         //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                       //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                       //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                       //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                      //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                      //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                         //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                       //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                      //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                      //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                        //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                      //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                       //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                      //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                     //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                      //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                     //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                      //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                     //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                     //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                         //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                       //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                       //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                       //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                      //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                      //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                          //                                                  clk_0_clk.clk
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),               // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),               //              onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.onchip_memory2_0_s1_address                                      (mm_interconnect_1_onchip_memory2_0_s1_address),    //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_1_onchip_memory2_0_s1_write),      //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_1_onchip_memory2_0_s1_clken)       //                                                           .clken
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                    //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                  //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                   //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                  //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                 //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                  //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                 //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                  //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                 //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                 //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                     //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                   //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                   //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                   //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                  //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                  //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                     //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                   //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                  //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                  //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                    //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                  //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                   //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                  //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                 //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                  //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                 //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                  //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                 //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                 //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                     //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                   //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                   //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                   //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                  //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                  //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                         //                                                     clk_0_clk.clk
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),              //              fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),              // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_reset_reset_bridge_in_reset_reset                      (rst_controller_001_reset_out_reset),              //                      lw_mm_bridge_reset_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                                     (fpga_only_master_master_address),                 //                                       fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                                 (fpga_only_master_master_waitrequest),             //                                                              .waitrequest
		.fpga_only_master_master_byteenable                                  (fpga_only_master_master_byteenable),              //                                                              .byteenable
		.fpga_only_master_master_read                                        (fpga_only_master_master_read),                    //                                                              .read
		.fpga_only_master_master_readdata                                    (fpga_only_master_master_readdata),                //                                                              .readdata
		.fpga_only_master_master_readdatavalid                               (fpga_only_master_master_readdatavalid),           //                                                              .readdatavalid
		.fpga_only_master_master_write                                       (fpga_only_master_master_write),                   //                                                              .write
		.fpga_only_master_master_writedata                                   (fpga_only_master_master_writedata),               //                                                              .writedata
		.lw_mm_bridge_s0_address                                             (mm_interconnect_2_lw_mm_bridge_s0_address),       //                                               lw_mm_bridge_s0.address
		.lw_mm_bridge_s0_write                                               (mm_interconnect_2_lw_mm_bridge_s0_write),         //                                                              .write
		.lw_mm_bridge_s0_read                                                (mm_interconnect_2_lw_mm_bridge_s0_read),          //                                                              .read
		.lw_mm_bridge_s0_readdata                                            (mm_interconnect_2_lw_mm_bridge_s0_readdata),      //                                                              .readdata
		.lw_mm_bridge_s0_writedata                                           (mm_interconnect_2_lw_mm_bridge_s0_writedata),     //                                                              .writedata
		.lw_mm_bridge_s0_burstcount                                          (mm_interconnect_2_lw_mm_bridge_s0_burstcount),    //                                                              .burstcount
		.lw_mm_bridge_s0_byteenable                                          (mm_interconnect_2_lw_mm_bridge_s0_byteenable),    //                                                              .byteenable
		.lw_mm_bridge_s0_readdatavalid                                       (mm_interconnect_2_lw_mm_bridge_s0_readdatavalid), //                                                              .readdatavalid
		.lw_mm_bridge_s0_waitrequest                                         (mm_interconnect_2_lw_mm_bridge_s0_waitrequest),   //                                                              .waitrequest
		.lw_mm_bridge_s0_debugaccess                                         (mm_interconnect_2_lw_mm_bridge_s0_debugaccess)    //                                                              .debugaccess
	);

	soc_system_mm_interconnect_3 mm_interconnect_3 (
		.clk_0_clk_clk                                           (clk_clk),                                                   //                                         clk_0_clk.clk
		.hps_0_h2f_user0_clock_clk                               (hps_0_h2f_user0_clock_clk),                                 //                             hps_0_h2f_user0_clock.clk
		.fft_sub_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                            //               fft_sub_reset_reset_bridge_in_reset.reset
		.fft_sub_s0_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // fft_sub_s0_translator_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_reset_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                        //          lw_mm_bridge_reset_reset_bridge_in_reset.reset
		.lw_mm_bridge_m0_address                                 (lw_mm_bridge_m0_address),                                   //                                   lw_mm_bridge_m0.address
		.lw_mm_bridge_m0_waitrequest                             (lw_mm_bridge_m0_waitrequest),                               //                                                  .waitrequest
		.lw_mm_bridge_m0_burstcount                              (lw_mm_bridge_m0_burstcount),                                //                                                  .burstcount
		.lw_mm_bridge_m0_byteenable                              (lw_mm_bridge_m0_byteenable),                                //                                                  .byteenable
		.lw_mm_bridge_m0_read                                    (lw_mm_bridge_m0_read),                                      //                                                  .read
		.lw_mm_bridge_m0_readdata                                (lw_mm_bridge_m0_readdata),                                  //                                                  .readdata
		.lw_mm_bridge_m0_readdatavalid                           (lw_mm_bridge_m0_readdatavalid),                             //                                                  .readdatavalid
		.lw_mm_bridge_m0_write                                   (lw_mm_bridge_m0_write),                                     //                                                  .write
		.lw_mm_bridge_m0_writedata                               (lw_mm_bridge_m0_writedata),                                 //                                                  .writedata
		.lw_mm_bridge_m0_debugaccess                             (lw_mm_bridge_m0_debugaccess),                               //                                                  .debugaccess
		.button_pio_s1_address                                   (mm_interconnect_3_button_pio_s1_address),                   //                                     button_pio_s1.address
		.button_pio_s1_write                                     (mm_interconnect_3_button_pio_s1_write),                     //                                                  .write
		.button_pio_s1_readdata                                  (mm_interconnect_3_button_pio_s1_readdata),                  //                                                  .readdata
		.button_pio_s1_writedata                                 (mm_interconnect_3_button_pio_s1_writedata),                 //                                                  .writedata
		.button_pio_s1_chipselect                                (mm_interconnect_3_button_pio_s1_chipselect),                //                                                  .chipselect
		.chip_id_read_mm_0_s0_read                               (mm_interconnect_3_chip_id_read_mm_0_s0_read),               //                              chip_id_read_mm_0_s0.read
		.chip_id_read_mm_0_s0_readdata                           (mm_interconnect_3_chip_id_read_mm_0_s0_readdata),           //                                                  .readdata
		.dipsw_pio_s1_address                                    (mm_interconnect_3_dipsw_pio_s1_address),                    //                                      dipsw_pio_s1.address
		.dipsw_pio_s1_write                                      (mm_interconnect_3_dipsw_pio_s1_write),                      //                                                  .write
		.dipsw_pio_s1_readdata                                   (mm_interconnect_3_dipsw_pio_s1_readdata),                   //                                                  .readdata
		.dipsw_pio_s1_writedata                                  (mm_interconnect_3_dipsw_pio_s1_writedata),                  //                                                  .writedata
		.dipsw_pio_s1_chipselect                                 (mm_interconnect_3_dipsw_pio_s1_chipselect),                 //                                                  .chipselect
		.fft_sub_s0_address                                      (mm_interconnect_3_fft_sub_s0_address),                      //                                        fft_sub_s0.address
		.fft_sub_s0_write                                        (mm_interconnect_3_fft_sub_s0_write),                        //                                                  .write
		.fft_sub_s0_read                                         (mm_interconnect_3_fft_sub_s0_read),                         //                                                  .read
		.fft_sub_s0_readdata                                     (mm_interconnect_3_fft_sub_s0_readdata),                     //                                                  .readdata
		.fft_sub_s0_writedata                                    (mm_interconnect_3_fft_sub_s0_writedata),                    //                                                  .writedata
		.fft_sub_s0_burstcount                                   (mm_interconnect_3_fft_sub_s0_burstcount),                   //                                                  .burstcount
		.fft_sub_s0_byteenable                                   (mm_interconnect_3_fft_sub_s0_byteenable),                   //                                                  .byteenable
		.fft_sub_s0_readdatavalid                                (mm_interconnect_3_fft_sub_s0_readdatavalid),                //                                                  .readdatavalid
		.fft_sub_s0_waitrequest                                  (mm_interconnect_3_fft_sub_s0_waitrequest),                  //                                                  .waitrequest
		.fft_sub_s0_debugaccess                                  (mm_interconnect_3_fft_sub_s0_debugaccess),                  //                                                  .debugaccess
		.intr_capturer_0_avalon_slave_0_address                  (mm_interconnect_3_intr_capturer_0_avalon_slave_0_address),  //                    intr_capturer_0_avalon_slave_0.address
		.intr_capturer_0_avalon_slave_0_read                     (mm_interconnect_3_intr_capturer_0_avalon_slave_0_read),     //                                                  .read
		.intr_capturer_0_avalon_slave_0_readdata                 (mm_interconnect_3_intr_capturer_0_avalon_slave_0_readdata), //                                                  .readdata
		.jtag_uart_avalon_jtag_slave_address                     (mm_interconnect_3_jtag_uart_avalon_jtag_slave_address),     //                       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                       (mm_interconnect_3_jtag_uart_avalon_jtag_slave_write),       //                                                  .write
		.jtag_uart_avalon_jtag_slave_read                        (mm_interconnect_3_jtag_uart_avalon_jtag_slave_read),        //                                                  .read
		.jtag_uart_avalon_jtag_slave_readdata                    (mm_interconnect_3_jtag_uart_avalon_jtag_slave_readdata),    //                                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata                   (mm_interconnect_3_jtag_uart_avalon_jtag_slave_writedata),   //                                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                 (mm_interconnect_3_jtag_uart_avalon_jtag_slave_waitrequest), //                                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                  (mm_interconnect_3_jtag_uart_avalon_jtag_slave_chipselect),  //                                                  .chipselect
		.led_pio_s1_address                                      (mm_interconnect_3_led_pio_s1_address),                      //                                        led_pio_s1.address
		.led_pio_s1_write                                        (mm_interconnect_3_led_pio_s1_write),                        //                                                  .write
		.led_pio_s1_readdata                                     (mm_interconnect_3_led_pio_s1_readdata),                     //                                                  .readdata
		.led_pio_s1_writedata                                    (mm_interconnect_3_led_pio_s1_writedata),                    //                                                  .writedata
		.led_pio_s1_chipselect                                   (mm_interconnect_3_led_pio_s1_chipselect),                   //                                                  .chipselect
		.sysid_qsys_control_slave_address                        (mm_interconnect_3_sysid_qsys_control_slave_address),        //                          sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                       (mm_interconnect_3_sysid_qsys_control_slave_readdata)        //                                                  .readdata
	);

	soc_system_mm_interconnect_5 mm_interconnect_5 (
		.hps_0_f2h_sdram0_data_awid                                              (mm_interconnect_5_hps_0_f2h_sdram0_data_awid),    //                                             hps_0_f2h_sdram0_data.awid
		.hps_0_f2h_sdram0_data_awaddr                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_awaddr),  //                                                                  .awaddr
		.hps_0_f2h_sdram0_data_awlen                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_awlen),   //                                                                  .awlen
		.hps_0_f2h_sdram0_data_awsize                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_awsize),  //                                                                  .awsize
		.hps_0_f2h_sdram0_data_awburst                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_awburst), //                                                                  .awburst
		.hps_0_f2h_sdram0_data_awlock                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_awlock),  //                                                                  .awlock
		.hps_0_f2h_sdram0_data_awcache                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_awcache), //                                                                  .awcache
		.hps_0_f2h_sdram0_data_awprot                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_awprot),  //                                                                  .awprot
		.hps_0_f2h_sdram0_data_awvalid                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_awvalid), //                                                                  .awvalid
		.hps_0_f2h_sdram0_data_awready                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_awready), //                                                                  .awready
		.hps_0_f2h_sdram0_data_wid                                               (mm_interconnect_5_hps_0_f2h_sdram0_data_wid),     //                                                                  .wid
		.hps_0_f2h_sdram0_data_wdata                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_wdata),   //                                                                  .wdata
		.hps_0_f2h_sdram0_data_wstrb                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_wstrb),   //                                                                  .wstrb
		.hps_0_f2h_sdram0_data_wlast                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_wlast),   //                                                                  .wlast
		.hps_0_f2h_sdram0_data_wvalid                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_wvalid),  //                                                                  .wvalid
		.hps_0_f2h_sdram0_data_wready                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_wready),  //                                                                  .wready
		.hps_0_f2h_sdram0_data_bid                                               (mm_interconnect_5_hps_0_f2h_sdram0_data_bid),     //                                                                  .bid
		.hps_0_f2h_sdram0_data_bresp                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_bresp),   //                                                                  .bresp
		.hps_0_f2h_sdram0_data_bvalid                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_bvalid),  //                                                                  .bvalid
		.hps_0_f2h_sdram0_data_bready                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_bready),  //                                                                  .bready
		.hps_0_f2h_sdram0_data_arid                                              (mm_interconnect_5_hps_0_f2h_sdram0_data_arid),    //                                                                  .arid
		.hps_0_f2h_sdram0_data_araddr                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_araddr),  //                                                                  .araddr
		.hps_0_f2h_sdram0_data_arlen                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_arlen),   //                                                                  .arlen
		.hps_0_f2h_sdram0_data_arsize                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_arsize),  //                                                                  .arsize
		.hps_0_f2h_sdram0_data_arburst                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_arburst), //                                                                  .arburst
		.hps_0_f2h_sdram0_data_arlock                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_arlock),  //                                                                  .arlock
		.hps_0_f2h_sdram0_data_arcache                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_arcache), //                                                                  .arcache
		.hps_0_f2h_sdram0_data_arprot                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_arprot),  //                                                                  .arprot
		.hps_0_f2h_sdram0_data_arvalid                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_arvalid), //                                                                  .arvalid
		.hps_0_f2h_sdram0_data_arready                                           (mm_interconnect_5_hps_0_f2h_sdram0_data_arready), //                                                                  .arready
		.hps_0_f2h_sdram0_data_rid                                               (mm_interconnect_5_hps_0_f2h_sdram0_data_rid),     //                                                                  .rid
		.hps_0_f2h_sdram0_data_rdata                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_rdata),   //                                                                  .rdata
		.hps_0_f2h_sdram0_data_rresp                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_rresp),   //                                                                  .rresp
		.hps_0_f2h_sdram0_data_rlast                                             (mm_interconnect_5_hps_0_f2h_sdram0_data_rlast),   //                                                                  .rlast
		.hps_0_f2h_sdram0_data_rvalid                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_rvalid),  //                                                                  .rvalid
		.hps_0_f2h_sdram0_data_rready                                            (mm_interconnect_5_hps_0_f2h_sdram0_data_rready),  //                                                                  .rready
		.clk_0_clk_clk                                                           (clk_clk),                                         //                                                         clk_0_clk.clk
		.f2sdram_only_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),              //               f2sdram_only_master_clk_reset_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),              // f2sdram_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_sdram0_data_agent_reset_sink_reset_bridge_in_reset_reset      (rst_controller_002_reset_out_reset),              //      hps_0_f2h_sdram0_data_agent_reset_sink_reset_bridge_in_reset.reset
		.f2sdram_only_master_master_address                                      (f2sdram_only_master_master_address),              //                                        f2sdram_only_master_master.address
		.f2sdram_only_master_master_waitrequest                                  (f2sdram_only_master_master_waitrequest),          //                                                                  .waitrequest
		.f2sdram_only_master_master_byteenable                                   (f2sdram_only_master_master_byteenable),           //                                                                  .byteenable
		.f2sdram_only_master_master_read                                         (f2sdram_only_master_master_read),                 //                                                                  .read
		.f2sdram_only_master_master_readdata                                     (f2sdram_only_master_master_readdata),             //                                                                  .readdata
		.f2sdram_only_master_master_readdatavalid                                (f2sdram_only_master_master_readdatavalid),        //                                                                  .readdatavalid
		.f2sdram_only_master_master_write                                        (f2sdram_only_master_master_write),                //                                                                  .write
		.f2sdram_only_master_master_writedata                                    (f2sdram_only_master_master_writedata)             //                                                                  .writedata
	);

	soc_system_mm_interconnect_6 mm_interconnect_6 (
		.hps_0_h2f_user0_clock_clk                        (hps_0_h2f_user0_clock_clk),                                     //                      hps_0_h2f_user0_clock.clk
		.fft_ddr_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // fft_ddr_bridge_reset_reset_bridge_in_reset.reset
		.fft_sub_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                //        fft_sub_reset_reset_bridge_in_reset.reset
		.fft_sub_to_ddr_address                           (fft_sub_to_ddr_address),                                        //                             fft_sub_to_ddr.address
		.fft_sub_to_ddr_waitrequest                       (fft_sub_to_ddr_waitrequest),                                    //                                           .waitrequest
		.fft_sub_to_ddr_burstcount                        (fft_sub_to_ddr_burstcount),                                     //                                           .burstcount
		.fft_sub_to_ddr_byteenable                        (fft_sub_to_ddr_byteenable),                                     //                                           .byteenable
		.fft_sub_to_ddr_read                              (fft_sub_to_ddr_read),                                           //                                           .read
		.fft_sub_to_ddr_readdata                          (fft_sub_to_ddr_readdata),                                       //                                           .readdata
		.fft_sub_to_ddr_readdatavalid                     (fft_sub_to_ddr_readdatavalid),                                  //                                           .readdatavalid
		.fft_sub_to_ddr_write                             (fft_sub_to_ddr_write),                                          //                                           .write
		.fft_sub_to_ddr_writedata                         (fft_sub_to_ddr_writedata),                                      //                                           .writedata
		.fft_sub_to_ddr_debugaccess                       (fft_sub_to_ddr_debugaccess),                                    //                                           .debugaccess
		.fft_ddr_bridge_windowed_slave_address            (mm_interconnect_6_fft_ddr_bridge_windowed_slave_address),       //              fft_ddr_bridge_windowed_slave.address
		.fft_ddr_bridge_windowed_slave_write              (mm_interconnect_6_fft_ddr_bridge_windowed_slave_write),         //                                           .write
		.fft_ddr_bridge_windowed_slave_read               (mm_interconnect_6_fft_ddr_bridge_windowed_slave_read),          //                                           .read
		.fft_ddr_bridge_windowed_slave_readdata           (mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdata),      //                                           .readdata
		.fft_ddr_bridge_windowed_slave_writedata          (mm_interconnect_6_fft_ddr_bridge_windowed_slave_writedata),     //                                           .writedata
		.fft_ddr_bridge_windowed_slave_burstcount         (mm_interconnect_6_fft_ddr_bridge_windowed_slave_burstcount),    //                                           .burstcount
		.fft_ddr_bridge_windowed_slave_byteenable         (mm_interconnect_6_fft_ddr_bridge_windowed_slave_byteenable),    //                                           .byteenable
		.fft_ddr_bridge_windowed_slave_readdatavalid      (mm_interconnect_6_fft_ddr_bridge_windowed_slave_readdatavalid), //                                           .readdatavalid
		.fft_ddr_bridge_windowed_slave_waitrequest        (mm_interconnect_6_fft_ddr_bridge_windowed_slave_waitrequest)    //                                           .waitrequest
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq), // receiver5.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_002 (
		.clk           (clk_clk),                                //       clk.clk
		.reset         (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),               // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),               // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),               // receiver2.irq
		.receiver3_irq (irq_mapper_002_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_002_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_002_receiver5_irq),           // receiver5.irq
		.sender_irq    (intr_capturer_0_interrupt_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (hps_0_h2f_user0_clock_clk),          //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_mapper_receiver3_irq),           //           receiver.irq
		.sender_irq     (irq_mapper_002_receiver3_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (hps_0_h2f_user0_clock_clk),          //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_mapper_receiver4_irq),           //           receiver.irq
		.sender_irq     (irq_mapper_002_receiver4_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (hps_0_h2f_user0_clock_clk),          //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_mapper_receiver5_irq),           //           receiver.irq
		.sender_irq     (irq_mapper_002_receiver5_irq)        //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (hps_0_h2f_user0_clock_clk),      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
