// soc_system_fft_sub.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module soc_system_fft_sub (
		input  wire        clk_clk,                    //                    clk.clk
		input  wire        reset_reset_n,              //                  reset.reset_n
		output wire        s0_waitrequest,             //                     s0.waitrequest
		output wire [31:0] s0_readdata,                //                       .readdata
		output wire        s0_readdatavalid,           //                       .readdatavalid
		input  wire [0:0]  s0_burstcount,              //                       .burstcount
		input  wire [31:0] s0_writedata,               //                       .writedata
		input  wire [18:0] s0_address,                 //                       .address
		input  wire        s0_write,                   //                       .write
		input  wire        s0_read,                    //                       .read
		input  wire [3:0]  s0_byteenable,              //                       .byteenable
		input  wire        s0_debugaccess,             //                       .debugaccess
		output wire        sgdma_from_fft_csr_irq_irq, // sgdma_from_fft_csr_irq.irq
		output wire        sgdma_from_ram_csr_irq_irq, // sgdma_from_ram_csr_irq.irq
		output wire        sgdma_to_fft_csr_irq_irq,   //   sgdma_to_fft_csr_irq.irq
		input  wire        to_ddr_waitrequest,         //                 to_ddr.waitrequest
		input  wire [63:0] to_ddr_readdata,            //                       .readdata
		input  wire        to_ddr_readdatavalid,       //                       .readdatavalid
		output wire [5:0]  to_ddr_burstcount,          //                       .burstcount
		output wire [63:0] to_ddr_writedata,           //                       .writedata
		output wire [29:0] to_ddr_address,             //                       .address
		output wire        to_ddr_write,               //                       .write
		output wire        to_ddr_read,                //                       .read
		output wire [7:0]  to_ddr_byteenable,          //                       .byteenable
		output wire        to_ddr_debugaccess          //                       .debugaccess
	);

	wire          fft_stadapter_0_out0_valid;                                    // FFT_STadapter_0:aso_out0_valid -> sgdma_from_fft:st_sink_valid
	wire   [63:0] fft_stadapter_0_out0_data;                                     // FFT_STadapter_0:aso_out0_data -> sgdma_from_fft:st_sink_data
	wire          fft_stadapter_0_out0_ready;                                    // sgdma_from_fft:st_sink_ready -> FFT_STadapter_0:aso_out0_ready
	wire          fft_stadapter_0_out0_startofpacket;                            // FFT_STadapter_0:aso_out0_startofpacket -> sgdma_from_fft:st_sink_startofpacket
	wire          fft_stadapter_0_out0_endofpacket;                              // FFT_STadapter_0:aso_out0_endofpacket -> sgdma_from_fft:st_sink_endofpacket
	wire    [1:0] fft_stadapter_0_out0_error;                                    // FFT_STadapter_0:aso_out0_error -> sgdma_from_fft:st_sink_error
	wire    [2:0] fft_stadapter_0_out0_empty;                                    // FFT_STadapter_0:aso_out0_empty -> sgdma_from_fft:st_sink_empty
	wire          fft_ii_0_source_valid;                                         // fft_ii_0:source_valid -> FFT_STadapter_0:asi_fromfft_valid
	wire   [61:0] fft_ii_0_source_data;                                          // fft_ii_0:source_data -> FFT_STadapter_0:asi_fromfft_data
	wire          fft_ii_0_source_ready;                                         // FFT_STadapter_0:asi_fromfft_ready -> fft_ii_0:source_ready
	wire          fft_ii_0_source_startofpacket;                                 // fft_ii_0:source_sop -> FFT_STadapter_0:asi_fromfft_startofpacket
	wire    [1:0] fft_ii_0_source_error;                                         // fft_ii_0:source_error -> FFT_STadapter_0:asi_fromfft_error
	wire          fft_ii_0_source_endofpacket;                                   // fft_ii_0:source_eop -> FFT_STadapter_0:asi_fromfft_endofpacket
	wire          sgdma_to_fft_st_source_valid;                                  // sgdma_to_fft:st_source_valid -> FFT_STadapter_0:asi_in0_valid
	wire   [31:0] sgdma_to_fft_st_source_data;                                   // sgdma_to_fft:st_source_data -> FFT_STadapter_0:asi_in0_data
	wire          sgdma_to_fft_st_source_ready;                                  // FFT_STadapter_0:asi_in0_ready -> sgdma_to_fft:st_source_ready
	wire          sgdma_to_fft_st_source_startofpacket;                          // sgdma_to_fft:st_source_startofpacket -> FFT_STadapter_0:asi_in0_startofpacket
	wire          sgdma_to_fft_st_source_endofpacket;                            // sgdma_to_fft:st_source_endofpacket -> FFT_STadapter_0:asi_in0_endofpacket
	wire    [1:0] sgdma_to_fft_st_source_error;                                  // sgdma_to_fft:st_source_error -> FFT_STadapter_0:asi_in0_error
	wire    [1:0] sgdma_to_fft_st_source_empty;                                  // sgdma_to_fft:st_source_empty -> FFT_STadapter_0:asi_in0_empty
	wire          fft_stadapter_0_tofft_valid;                                   // FFT_STadapter_0:aso_tofft_valid -> fft_ii_0:sink_valid
	wire   [46:0] fft_stadapter_0_tofft_data;                                    // FFT_STadapter_0:aso_tofft_data -> fft_ii_0:sink_data
	wire          fft_stadapter_0_tofft_ready;                                   // fft_ii_0:sink_ready -> FFT_STadapter_0:aso_tofft_ready
	wire          fft_stadapter_0_tofft_startofpacket;                           // FFT_STadapter_0:aso_tofft_startofpacket -> fft_ii_0:sink_sop
	wire          fft_stadapter_0_tofft_endofpacket;                             // FFT_STadapter_0:aso_tofft_endofpacket -> fft_ii_0:sink_eop
	wire    [1:0] fft_stadapter_0_tofft_error;                                   // FFT_STadapter_0:aso_tofft_error -> fft_ii_0:sink_error
	wire          mm_bridge_0_m0_waitrequest;                                    // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire   [31:0] mm_bridge_0_m0_readdata;                                       // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire          mm_bridge_0_m0_debugaccess;                                    // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [18:0] mm_bridge_0_m0_address;                                        // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire          mm_bridge_0_m0_read;                                           // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire    [3:0] mm_bridge_0_m0_byteenable;                                     // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire          mm_bridge_0_m0_readdatavalid;                                  // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire   [31:0] mm_bridge_0_m0_writedata;                                      // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire          mm_bridge_0_m0_write;                                          // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire    [0:0] mm_bridge_0_m0_burstcount;                                     // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire   [31:0] sgdma_to_fft_mm_read_readdata;                                 // mm_interconnect_0:sgdma_to_fft_mm_read_readdata -> sgdma_to_fft:mm_read_readdata
	wire          sgdma_to_fft_mm_read_waitrequest;                              // mm_interconnect_0:sgdma_to_fft_mm_read_waitrequest -> sgdma_to_fft:mm_read_waitrequest
	wire   [30:0] sgdma_to_fft_mm_read_address;                                  // sgdma_to_fft:mm_read_address -> mm_interconnect_0:sgdma_to_fft_mm_read_address
	wire          sgdma_to_fft_mm_read_read;                                     // sgdma_to_fft:mm_read_read -> mm_interconnect_0:sgdma_to_fft_mm_read_read
	wire    [3:0] sgdma_to_fft_mm_read_byteenable;                               // sgdma_to_fft:mm_read_byteenable -> mm_interconnect_0:sgdma_to_fft_mm_read_byteenable
	wire          sgdma_to_fft_mm_read_readdatavalid;                            // mm_interconnect_0:sgdma_to_fft_mm_read_readdatavalid -> sgdma_to_fft:mm_read_readdatavalid
	wire    [6:0] sgdma_to_fft_mm_read_burstcount;                               // sgdma_to_fft:mm_read_burstcount -> mm_interconnect_0:sgdma_to_fft_mm_read_burstcount
	wire   [63:0] sgdma_from_ram_mm_read_readdata;                               // mm_interconnect_0:sgdma_from_ram_mm_read_readdata -> sgdma_from_ram:mm_read_readdata
	wire          sgdma_from_ram_mm_read_waitrequest;                            // mm_interconnect_0:sgdma_from_ram_mm_read_waitrequest -> sgdma_from_ram:mm_read_waitrequest
	wire   [18:0] sgdma_from_ram_mm_read_address;                                // sgdma_from_ram:mm_read_address -> mm_interconnect_0:sgdma_from_ram_mm_read_address
	wire          sgdma_from_ram_mm_read_read;                                   // sgdma_from_ram:mm_read_read -> mm_interconnect_0:sgdma_from_ram_mm_read_read
	wire    [7:0] sgdma_from_ram_mm_read_byteenable;                             // sgdma_from_ram:mm_read_byteenable -> mm_interconnect_0:sgdma_from_ram_mm_read_byteenable
	wire          sgdma_from_ram_mm_read_readdatavalid;                          // mm_interconnect_0:sgdma_from_ram_mm_read_readdatavalid -> sgdma_from_ram:mm_read_readdatavalid
	wire    [5:0] sgdma_from_ram_mm_read_burstcount;                             // sgdma_from_ram:mm_read_burstcount -> mm_interconnect_0:sgdma_from_ram_mm_read_burstcount
	wire          sgdma_from_fft_mm_write_waitrequest;                           // mm_interconnect_0:sgdma_from_fft_mm_write_waitrequest -> sgdma_from_fft:mm_write_waitrequest
	wire   [30:0] sgdma_from_fft_mm_write_address;                               // sgdma_from_fft:mm_write_address -> mm_interconnect_0:sgdma_from_fft_mm_write_address
	wire    [7:0] sgdma_from_fft_mm_write_byteenable;                            // sgdma_from_fft:mm_write_byteenable -> mm_interconnect_0:sgdma_from_fft_mm_write_byteenable
	wire          sgdma_from_fft_mm_write_write;                                 // sgdma_from_fft:mm_write_write -> mm_interconnect_0:sgdma_from_fft_mm_write_write
	wire   [63:0] sgdma_from_fft_mm_write_writedata;                             // sgdma_from_fft:mm_write_writedata -> mm_interconnect_0:sgdma_from_fft_mm_write_writedata
	wire    [5:0] sgdma_from_fft_mm_write_burstcount;                            // sgdma_from_fft:mm_write_burstcount -> mm_interconnect_0:sgdma_from_fft_mm_write_burstcount
	wire          sgdma_from_ram_mm_write_waitrequest;                           // mm_interconnect_0:sgdma_from_ram_mm_write_waitrequest -> sgdma_from_ram:mm_write_waitrequest
	wire   [30:0] sgdma_from_ram_mm_write_address;                               // sgdma_from_ram:mm_write_address -> mm_interconnect_0:sgdma_from_ram_mm_write_address
	wire    [7:0] sgdma_from_ram_mm_write_byteenable;                            // sgdma_from_ram:mm_write_byteenable -> mm_interconnect_0:sgdma_from_ram_mm_write_byteenable
	wire          sgdma_from_ram_mm_write_write;                                 // sgdma_from_ram:mm_write_write -> mm_interconnect_0:sgdma_from_ram_mm_write_write
	wire   [63:0] sgdma_from_ram_mm_write_writedata;                             // sgdma_from_ram:mm_write_writedata -> mm_interconnect_0:sgdma_from_ram_mm_write_writedata
	wire    [5:0] sgdma_from_ram_mm_write_burstcount;                            // sgdma_from_ram:mm_write_burstcount -> mm_interconnect_0:sgdma_from_ram_mm_write_burstcount
	wire   [31:0] mm_interconnect_0_sgdma_from_fft_csr_readdata;                 // sgdma_from_fft:csr_readdata -> mm_interconnect_0:sgdma_from_fft_csr_readdata
	wire    [2:0] mm_interconnect_0_sgdma_from_fft_csr_address;                  // mm_interconnect_0:sgdma_from_fft_csr_address -> sgdma_from_fft:csr_address
	wire          mm_interconnect_0_sgdma_from_fft_csr_read;                     // mm_interconnect_0:sgdma_from_fft_csr_read -> sgdma_from_fft:csr_read
	wire    [3:0] mm_interconnect_0_sgdma_from_fft_csr_byteenable;               // mm_interconnect_0:sgdma_from_fft_csr_byteenable -> sgdma_from_fft:csr_byteenable
	wire          mm_interconnect_0_sgdma_from_fft_csr_write;                    // mm_interconnect_0:sgdma_from_fft_csr_write -> sgdma_from_fft:csr_write
	wire   [31:0] mm_interconnect_0_sgdma_from_fft_csr_writedata;                // mm_interconnect_0:sgdma_from_fft_csr_writedata -> sgdma_from_fft:csr_writedata
	wire   [31:0] mm_interconnect_0_sgdma_to_fft_csr_readdata;                   // sgdma_to_fft:csr_readdata -> mm_interconnect_0:sgdma_to_fft_csr_readdata
	wire    [2:0] mm_interconnect_0_sgdma_to_fft_csr_address;                    // mm_interconnect_0:sgdma_to_fft_csr_address -> sgdma_to_fft:csr_address
	wire          mm_interconnect_0_sgdma_to_fft_csr_read;                       // mm_interconnect_0:sgdma_to_fft_csr_read -> sgdma_to_fft:csr_read
	wire    [3:0] mm_interconnect_0_sgdma_to_fft_csr_byteenable;                 // mm_interconnect_0:sgdma_to_fft_csr_byteenable -> sgdma_to_fft:csr_byteenable
	wire          mm_interconnect_0_sgdma_to_fft_csr_write;                      // mm_interconnect_0:sgdma_to_fft_csr_write -> sgdma_to_fft:csr_write
	wire   [31:0] mm_interconnect_0_sgdma_to_fft_csr_writedata;                  // mm_interconnect_0:sgdma_to_fft_csr_writedata -> sgdma_to_fft:csr_writedata
	wire   [31:0] mm_interconnect_0_sgdma_from_ram_csr_readdata;                 // sgdma_from_ram:csr_readdata -> mm_interconnect_0:sgdma_from_ram_csr_readdata
	wire    [2:0] mm_interconnect_0_sgdma_from_ram_csr_address;                  // mm_interconnect_0:sgdma_from_ram_csr_address -> sgdma_from_ram:csr_address
	wire          mm_interconnect_0_sgdma_from_ram_csr_read;                     // mm_interconnect_0:sgdma_from_ram_csr_read -> sgdma_from_ram:csr_read
	wire    [3:0] mm_interconnect_0_sgdma_from_ram_csr_byteenable;               // mm_interconnect_0:sgdma_from_ram_csr_byteenable -> sgdma_from_ram:csr_byteenable
	wire          mm_interconnect_0_sgdma_from_ram_csr_write;                    // mm_interconnect_0:sgdma_from_ram_csr_write -> sgdma_from_ram:csr_write
	wire   [31:0] mm_interconnect_0_sgdma_from_ram_csr_writedata;                // mm_interconnect_0:sgdma_from_ram_csr_writedata -> sgdma_from_ram:csr_writedata
	wire          mm_interconnect_0_sgdma_from_fft_descriptor_slave_waitrequest; // sgdma_from_fft:descriptor_slave_waitrequest -> mm_interconnect_0:sgdma_from_fft_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_sgdma_from_fft_descriptor_slave_byteenable;  // mm_interconnect_0:sgdma_from_fft_descriptor_slave_byteenable -> sgdma_from_fft:descriptor_slave_byteenable
	wire          mm_interconnect_0_sgdma_from_fft_descriptor_slave_write;       // mm_interconnect_0:sgdma_from_fft_descriptor_slave_write -> sgdma_from_fft:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_sgdma_from_fft_descriptor_slave_writedata;   // mm_interconnect_0:sgdma_from_fft_descriptor_slave_writedata -> sgdma_from_fft:descriptor_slave_writedata
	wire          mm_interconnect_0_sgdma_to_fft_descriptor_slave_waitrequest;   // sgdma_to_fft:descriptor_slave_waitrequest -> mm_interconnect_0:sgdma_to_fft_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_sgdma_to_fft_descriptor_slave_byteenable;    // mm_interconnect_0:sgdma_to_fft_descriptor_slave_byteenable -> sgdma_to_fft:descriptor_slave_byteenable
	wire          mm_interconnect_0_sgdma_to_fft_descriptor_slave_write;         // mm_interconnect_0:sgdma_to_fft_descriptor_slave_write -> sgdma_to_fft:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_sgdma_to_fft_descriptor_slave_writedata;     // mm_interconnect_0:sgdma_to_fft_descriptor_slave_writedata -> sgdma_to_fft:descriptor_slave_writedata
	wire          mm_interconnect_0_sgdma_from_ram_descriptor_slave_waitrequest; // sgdma_from_ram:descriptor_slave_waitrequest -> mm_interconnect_0:sgdma_from_ram_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_sgdma_from_ram_descriptor_slave_byteenable;  // mm_interconnect_0:sgdma_from_ram_descriptor_slave_byteenable -> sgdma_from_ram:descriptor_slave_byteenable
	wire          mm_interconnect_0_sgdma_from_ram_descriptor_slave_write;       // mm_interconnect_0:sgdma_from_ram_descriptor_slave_write -> sgdma_from_ram:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_sgdma_from_ram_descriptor_slave_writedata;   // mm_interconnect_0:sgdma_from_ram_descriptor_slave_writedata -> sgdma_from_ram:descriptor_slave_writedata
	wire   [31:0] mm_interconnect_0_fft_stadapter_0_s0_readdata;                 // FFT_STadapter_0:avs_s0_readdata -> mm_interconnect_0:FFT_STadapter_0_s0_readdata
	wire    [1:0] mm_interconnect_0_fft_stadapter_0_s0_address;                  // mm_interconnect_0:FFT_STadapter_0_s0_address -> FFT_STadapter_0:avs_s0_address
	wire          mm_interconnect_0_fft_stadapter_0_s0_read;                     // mm_interconnect_0:FFT_STadapter_0_s0_read -> FFT_STadapter_0:avs_s0_read
	wire          mm_interconnect_0_fft_stadapter_0_s0_write;                    // mm_interconnect_0:FFT_STadapter_0_s0_write -> FFT_STadapter_0:avs_s0_write
	wire   [31:0] mm_interconnect_0_fft_stadapter_0_s0_writedata;                // mm_interconnect_0:FFT_STadapter_0_s0_writedata -> FFT_STadapter_0:avs_s0_writedata
	wire          mm_interconnect_0_data_s1_chipselect;                          // mm_interconnect_0:data_s1_chipselect -> data:chipselect
	wire   [63:0] mm_interconnect_0_data_s1_readdata;                            // data:readdata -> mm_interconnect_0:data_s1_readdata
	wire   [12:0] mm_interconnect_0_data_s1_address;                             // mm_interconnect_0:data_s1_address -> data:address
	wire    [7:0] mm_interconnect_0_data_s1_byteenable;                          // mm_interconnect_0:data_s1_byteenable -> data:byteenable
	wire          mm_interconnect_0_data_s1_write;                               // mm_interconnect_0:data_s1_write -> data:write
	wire   [63:0] mm_interconnect_0_data_s1_writedata;                           // mm_interconnect_0:data_s1_writedata -> data:writedata
	wire          mm_interconnect_0_data_s1_clken;                               // mm_interconnect_0:data_s1_clken -> data:clken
	wire   [63:0] mm_interconnect_0_ddr_s0_readdata;                             // DDR:s0_readdata -> mm_interconnect_0:DDR_s0_readdata
	wire          mm_interconnect_0_ddr_s0_waitrequest;                          // DDR:s0_waitrequest -> mm_interconnect_0:DDR_s0_waitrequest
	wire          mm_interconnect_0_ddr_s0_debugaccess;                          // mm_interconnect_0:DDR_s0_debugaccess -> DDR:s0_debugaccess
	wire   [29:0] mm_interconnect_0_ddr_s0_address;                              // mm_interconnect_0:DDR_s0_address -> DDR:s0_address
	wire          mm_interconnect_0_ddr_s0_read;                                 // mm_interconnect_0:DDR_s0_read -> DDR:s0_read
	wire    [7:0] mm_interconnect_0_ddr_s0_byteenable;                           // mm_interconnect_0:DDR_s0_byteenable -> DDR:s0_byteenable
	wire          mm_interconnect_0_ddr_s0_readdatavalid;                        // DDR:s0_readdatavalid -> mm_interconnect_0:DDR_s0_readdatavalid
	wire          mm_interconnect_0_ddr_s0_write;                                // mm_interconnect_0:DDR_s0_write -> DDR:s0_write
	wire   [63:0] mm_interconnect_0_ddr_s0_writedata;                            // mm_interconnect_0:DDR_s0_writedata -> DDR:s0_writedata
	wire    [5:0] mm_interconnect_0_ddr_s0_burstcount;                           // mm_interconnect_0:DDR_s0_burstcount -> DDR:s0_burstcount
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [DDR:reset, FFT_STadapter_0:reset, data:reset, fft_ii_0:reset_n, mm_bridge_0:reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sgdma_from_fft:reset_n_reset_n, sgdma_from_ram:reset_n_reset_n, sgdma_to_fft:reset_n_reset_n]
	wire          rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [data:reset_req, rst_translator:reset_req_in]
	wire   [23:0] fft_ii_0_source_imag;                                          // port fragment
	wire   [23:0] fft_ii_0_source_real;                                          // port fragment
	wire   [13:0] fft_ii_0_fftpts_out;                                           // port fragment

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (64),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (30),
		.BURSTCOUNT_WIDTH  (6),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) ddr (
		.clk              (clk_clk),                                //   clk.clk
		.reset            (rst_controller_reset_out_reset),         // reset.reset
		.s0_waitrequest   (mm_interconnect_0_ddr_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_ddr_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_ddr_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_ddr_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_ddr_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_ddr_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_ddr_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_ddr_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_ddr_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_ddr_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (to_ddr_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (to_ddr_readdata),                        //      .readdata
		.m0_readdatavalid (to_ddr_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (to_ddr_burstcount),                      //      .burstcount
		.m0_writedata     (to_ddr_writedata),                       //      .writedata
		.m0_address       (to_ddr_address),                         //      .address
		.m0_write         (to_ddr_write),                           //      .write
		.m0_read          (to_ddr_read),                            //      .read
		.m0_byteenable    (to_ddr_byteenable),                      //      .byteenable
		.m0_debugaccess   (to_ddr_debugaccess),                     //      .debugaccess
		.s0_response      (),                                       // (terminated)
		.m0_response      (2'b00)                                   // (terminated)
	);

	fft_adapter #(
		.FFT_IN_WIDTH  (16),
		.FFT_OUT_WIDTH (24),
		.SIZE_WIDTH    (14)
	) fft_stadapter_0 (
		.asi_in0_ready             (sgdma_to_fft_st_source_ready),                   //     in0.ready
		.asi_in0_valid             (sgdma_to_fft_st_source_valid),                   //        .valid
		.asi_in0_startofpacket     (sgdma_to_fft_st_source_startofpacket),           //        .startofpacket
		.asi_in0_endofpacket       (sgdma_to_fft_st_source_endofpacket),             //        .endofpacket
		.asi_in0_error             (sgdma_to_fft_st_source_error),                   //        .error
		.asi_in0_empty             (sgdma_to_fft_st_source_empty),                   //        .empty
		.asi_in0_data              (sgdma_to_fft_st_source_data),                    //        .data
		.clk                       (clk_clk),                                        //   clock.clk
		.reset                     (rst_controller_reset_out_reset),                 //   reset.reset
		.aso_out0_data             (fft_stadapter_0_out0_data),                      //    out0.data
		.aso_out0_ready            (fft_stadapter_0_out0_ready),                     //        .ready
		.aso_out0_valid            (fft_stadapter_0_out0_valid),                     //        .valid
		.aso_out0_startofpacket    (fft_stadapter_0_out0_startofpacket),             //        .startofpacket
		.aso_out0_endofpacket      (fft_stadapter_0_out0_endofpacket),               //        .endofpacket
		.aso_out0_error            (fft_stadapter_0_out0_error),                     //        .error
		.aso_out0_empty            (fft_stadapter_0_out0_empty),                     //        .empty
		.asi_fromfft_data          (fft_ii_0_source_data),                           // fromfft.data
		.asi_fromfft_ready         (fft_ii_0_source_ready),                          //        .ready
		.asi_fromfft_valid         (fft_ii_0_source_valid),                          //        .valid
		.asi_fromfft_startofpacket (fft_ii_0_source_startofpacket),                  //        .startofpacket
		.asi_fromfft_endofpacket   (fft_ii_0_source_endofpacket),                    //        .endofpacket
		.asi_fromfft_error         (fft_ii_0_source_error),                          //        .error
		.aso_tofft_data            (fft_stadapter_0_tofft_data),                     //   tofft.data
		.aso_tofft_ready           (fft_stadapter_0_tofft_ready),                    //        .ready
		.aso_tofft_valid           (fft_stadapter_0_tofft_valid),                    //        .valid
		.aso_tofft_startofpacket   (fft_stadapter_0_tofft_startofpacket),            //        .startofpacket
		.aso_tofft_endofpacket     (fft_stadapter_0_tofft_endofpacket),              //        .endofpacket
		.aso_tofft_error           (fft_stadapter_0_tofft_error),                    //        .error
		.avs_s0_address            (mm_interconnect_0_fft_stadapter_0_s0_address),   //      s0.address
		.avs_s0_read               (mm_interconnect_0_fft_stadapter_0_s0_read),      //        .read
		.avs_s0_readdata           (mm_interconnect_0_fft_stadapter_0_s0_readdata),  //        .readdata
		.avs_s0_write              (mm_interconnect_0_fft_stadapter_0_s0_write),     //        .write
		.avs_s0_writedata          (mm_interconnect_0_fft_stadapter_0_s0_writedata)  //        .writedata
	);

	soc_system_fft_sub_data data (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_data_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	soc_system_fft_sub_fft_ii_0 fft_ii_0 (
		.clk          (clk_clk),                             //    clk.clk
		.reset_n      (~rst_controller_reset_out_reset),     //    rst.reset_n
		.sink_valid   (fft_stadapter_0_tofft_valid),         //   sink.valid
		.sink_ready   (fft_stadapter_0_tofft_ready),         //       .ready
		.sink_error   (fft_stadapter_0_tofft_error),         //       .error
		.sink_sop     (fft_stadapter_0_tofft_startofpacket), //       .startofpacket
		.sink_eop     (fft_stadapter_0_tofft_endofpacket),   //       .endofpacket
		.sink_real    (fft_stadapter_0_tofft_data[46:31]),   //       .data
		.sink_imag    (fft_stadapter_0_tofft_data[30:15]),   //       .data
		.fftpts_in    (fft_stadapter_0_tofft_data[14:1]),    //       .data
		.inverse      (fft_stadapter_0_tofft_data[0]),       //       .data
		.source_valid (fft_ii_0_source_valid),               // source.valid
		.source_ready (fft_ii_0_source_ready),               //       .ready
		.source_error (fft_ii_0_source_error),               //       .error
		.source_sop   (fft_ii_0_source_startofpacket),       //       .startofpacket
		.source_eop   (fft_ii_0_source_endofpacket),         //       .endofpacket
		.source_real  (fft_ii_0_source_real[23:0]),          //       .data
		.source_imag  (fft_ii_0_source_imag[23:0]),          //       .data
		.fftpts_out   (fft_ii_0_fftpts_out[13:0])            //       .data
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (19),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                        //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (s0_waitrequest),                 //    s0.waitrequest
		.s0_readdata      (s0_readdata),                    //      .readdata
		.s0_readdatavalid (s0_readdatavalid),               //      .readdatavalid
		.s0_burstcount    (s0_burstcount),                  //      .burstcount
		.s0_writedata     (s0_writedata),                   //      .writedata
		.s0_address       (s0_address),                     //      .address
		.s0_write         (s0_write),                       //      .write
		.s0_read          (s0_read),                        //      .read
		.s0_byteenable    (s0_byteenable),                  //      .byteenable
		.s0_debugaccess   (s0_debugaccess),                 //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),         //      .address
		.m0_write         (mm_bridge_0_m0_write),           //      .write
		.m0_read          (mm_bridge_0_m0_read),            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess),     //      .debugaccess
		.s0_response      (),                               // (terminated)
		.m0_response      (2'b00)                           // (terminated)
	);

	soc_system_fft_sub_sgdma_from_fft sgdma_from_fft (
		.mm_write_address             (sgdma_from_fft_mm_write_address),                               //         mm_write.address
		.mm_write_write               (sgdma_from_fft_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (sgdma_from_fft_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (sgdma_from_fft_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (sgdma_from_fft_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (sgdma_from_fft_mm_write_burstcount),                            //                 .burstcount
		.clock_clk                    (clk_clk),                                                       //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                               //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_sgdma_from_fft_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_sgdma_from_fft_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_sgdma_from_fft_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_sgdma_from_fft_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_sgdma_from_fft_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_sgdma_from_fft_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_sgdma_from_fft_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_sgdma_from_fft_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_sgdma_from_fft_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_sgdma_from_fft_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (sgdma_from_fft_csr_irq_irq),                                    //          csr_irq.irq
		.st_sink_data                 (fft_stadapter_0_out0_data),                                     //          st_sink.data
		.st_sink_valid                (fft_stadapter_0_out0_valid),                                    //                 .valid
		.st_sink_ready                (fft_stadapter_0_out0_ready),                                    //                 .ready
		.st_sink_startofpacket        (fft_stadapter_0_out0_startofpacket),                            //                 .startofpacket
		.st_sink_endofpacket          (fft_stadapter_0_out0_endofpacket),                              //                 .endofpacket
		.st_sink_empty                (fft_stadapter_0_out0_empty),                                    //                 .empty
		.st_sink_error                (fft_stadapter_0_out0_error)                                     //                 .error
	);

	soc_system_fft_sub_sgdma_from_ram sgdma_from_ram (
		.mm_read_address              (sgdma_from_ram_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (sgdma_from_ram_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (sgdma_from_ram_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (sgdma_from_ram_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (sgdma_from_ram_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (sgdma_from_ram_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (sgdma_from_ram_mm_read_burstcount),                             //                 .burstcount
		.mm_write_address             (sgdma_from_ram_mm_write_address),                               //         mm_write.address
		.mm_write_write               (sgdma_from_ram_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (sgdma_from_ram_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (sgdma_from_ram_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (sgdma_from_ram_mm_write_waitrequest),                           //                 .waitrequest
		.mm_write_burstcount          (sgdma_from_ram_mm_write_burstcount),                            //                 .burstcount
		.clock_clk                    (clk_clk),                                                       //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                               //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_sgdma_from_ram_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_sgdma_from_ram_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_sgdma_from_ram_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_sgdma_from_ram_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_sgdma_from_ram_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_sgdma_from_ram_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_sgdma_from_ram_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_sgdma_from_ram_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_sgdma_from_ram_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_sgdma_from_ram_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (sgdma_from_ram_csr_irq_irq)                                     //          csr_irq.irq
	);

	soc_system_fft_sub_sgdma_to_fft sgdma_to_fft (
		.mm_read_address              (sgdma_to_fft_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (sgdma_to_fft_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (sgdma_to_fft_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (sgdma_to_fft_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (sgdma_to_fft_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (sgdma_to_fft_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_read_burstcount           (sgdma_to_fft_mm_read_burstcount),                             //                 .burstcount
		.clock_clk                    (clk_clk),                                                     //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                             //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_sgdma_to_fft_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_sgdma_to_fft_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_sgdma_to_fft_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_sgdma_to_fft_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_sgdma_to_fft_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_sgdma_to_fft_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_sgdma_to_fft_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_sgdma_to_fft_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_sgdma_to_fft_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_sgdma_to_fft_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (sgdma_to_fft_csr_irq_irq),                                    //          csr_irq.irq
		.st_source_data               (sgdma_to_fft_st_source_data),                                 //        st_source.data
		.st_source_valid              (sgdma_to_fft_st_source_valid),                                //                 .valid
		.st_source_ready              (sgdma_to_fft_st_source_ready),                                //                 .ready
		.st_source_startofpacket      (sgdma_to_fft_st_source_startofpacket),                        //                 .startofpacket
		.st_source_endofpacket        (sgdma_to_fft_st_source_endofpacket),                          //                 .endofpacket
		.st_source_empty              (sgdma_to_fft_st_source_empty),                                //                 .empty
		.st_source_error              (sgdma_to_fft_st_source_error)                                 //                 .error
	);

	soc_system_fft_sub_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                                       //                               clk_0_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                        //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                    //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                     //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                     //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                           //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                       //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                                  //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                          //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                      //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                    //                                        .debugaccess
		.sgdma_from_fft_mm_write_address               (sgdma_from_fft_mm_write_address),                               //                 sgdma_from_fft_mm_write.address
		.sgdma_from_fft_mm_write_waitrequest           (sgdma_from_fft_mm_write_waitrequest),                           //                                        .waitrequest
		.sgdma_from_fft_mm_write_burstcount            (sgdma_from_fft_mm_write_burstcount),                            //                                        .burstcount
		.sgdma_from_fft_mm_write_byteenable            (sgdma_from_fft_mm_write_byteenable),                            //                                        .byteenable
		.sgdma_from_fft_mm_write_write                 (sgdma_from_fft_mm_write_write),                                 //                                        .write
		.sgdma_from_fft_mm_write_writedata             (sgdma_from_fft_mm_write_writedata),                             //                                        .writedata
		.sgdma_from_ram_mm_read_address                (sgdma_from_ram_mm_read_address),                                //                  sgdma_from_ram_mm_read.address
		.sgdma_from_ram_mm_read_waitrequest            (sgdma_from_ram_mm_read_waitrequest),                            //                                        .waitrequest
		.sgdma_from_ram_mm_read_burstcount             (sgdma_from_ram_mm_read_burstcount),                             //                                        .burstcount
		.sgdma_from_ram_mm_read_byteenable             (sgdma_from_ram_mm_read_byteenable),                             //                                        .byteenable
		.sgdma_from_ram_mm_read_read                   (sgdma_from_ram_mm_read_read),                                   //                                        .read
		.sgdma_from_ram_mm_read_readdata               (sgdma_from_ram_mm_read_readdata),                               //                                        .readdata
		.sgdma_from_ram_mm_read_readdatavalid          (sgdma_from_ram_mm_read_readdatavalid),                          //                                        .readdatavalid
		.sgdma_from_ram_mm_write_address               (sgdma_from_ram_mm_write_address),                               //                 sgdma_from_ram_mm_write.address
		.sgdma_from_ram_mm_write_waitrequest           (sgdma_from_ram_mm_write_waitrequest),                           //                                        .waitrequest
		.sgdma_from_ram_mm_write_burstcount            (sgdma_from_ram_mm_write_burstcount),                            //                                        .burstcount
		.sgdma_from_ram_mm_write_byteenable            (sgdma_from_ram_mm_write_byteenable),                            //                                        .byteenable
		.sgdma_from_ram_mm_write_write                 (sgdma_from_ram_mm_write_write),                                 //                                        .write
		.sgdma_from_ram_mm_write_writedata             (sgdma_from_ram_mm_write_writedata),                             //                                        .writedata
		.sgdma_to_fft_mm_read_address                  (sgdma_to_fft_mm_read_address),                                  //                    sgdma_to_fft_mm_read.address
		.sgdma_to_fft_mm_read_waitrequest              (sgdma_to_fft_mm_read_waitrequest),                              //                                        .waitrequest
		.sgdma_to_fft_mm_read_burstcount               (sgdma_to_fft_mm_read_burstcount),                               //                                        .burstcount
		.sgdma_to_fft_mm_read_byteenable               (sgdma_to_fft_mm_read_byteenable),                               //                                        .byteenable
		.sgdma_to_fft_mm_read_read                     (sgdma_to_fft_mm_read_read),                                     //                                        .read
		.sgdma_to_fft_mm_read_readdata                 (sgdma_to_fft_mm_read_readdata),                                 //                                        .readdata
		.sgdma_to_fft_mm_read_readdatavalid            (sgdma_to_fft_mm_read_readdatavalid),                            //                                        .readdatavalid
		.data_s1_address                               (mm_interconnect_0_data_s1_address),                             //                                 data_s1.address
		.data_s1_write                                 (mm_interconnect_0_data_s1_write),                               //                                        .write
		.data_s1_readdata                              (mm_interconnect_0_data_s1_readdata),                            //                                        .readdata
		.data_s1_writedata                             (mm_interconnect_0_data_s1_writedata),                           //                                        .writedata
		.data_s1_byteenable                            (mm_interconnect_0_data_s1_byteenable),                          //                                        .byteenable
		.data_s1_chipselect                            (mm_interconnect_0_data_s1_chipselect),                          //                                        .chipselect
		.data_s1_clken                                 (mm_interconnect_0_data_s1_clken),                               //                                        .clken
		.DDR_s0_address                                (mm_interconnect_0_ddr_s0_address),                              //                                  DDR_s0.address
		.DDR_s0_write                                  (mm_interconnect_0_ddr_s0_write),                                //                                        .write
		.DDR_s0_read                                   (mm_interconnect_0_ddr_s0_read),                                 //                                        .read
		.DDR_s0_readdata                               (mm_interconnect_0_ddr_s0_readdata),                             //                                        .readdata
		.DDR_s0_writedata                              (mm_interconnect_0_ddr_s0_writedata),                            //                                        .writedata
		.DDR_s0_burstcount                             (mm_interconnect_0_ddr_s0_burstcount),                           //                                        .burstcount
		.DDR_s0_byteenable                             (mm_interconnect_0_ddr_s0_byteenable),                           //                                        .byteenable
		.DDR_s0_readdatavalid                          (mm_interconnect_0_ddr_s0_readdatavalid),                        //                                        .readdatavalid
		.DDR_s0_waitrequest                            (mm_interconnect_0_ddr_s0_waitrequest),                          //                                        .waitrequest
		.DDR_s0_debugaccess                            (mm_interconnect_0_ddr_s0_debugaccess),                          //                                        .debugaccess
		.FFT_STadapter_0_s0_address                    (mm_interconnect_0_fft_stadapter_0_s0_address),                  //                      FFT_STadapter_0_s0.address
		.FFT_STadapter_0_s0_write                      (mm_interconnect_0_fft_stadapter_0_s0_write),                    //                                        .write
		.FFT_STadapter_0_s0_read                       (mm_interconnect_0_fft_stadapter_0_s0_read),                     //                                        .read
		.FFT_STadapter_0_s0_readdata                   (mm_interconnect_0_fft_stadapter_0_s0_readdata),                 //                                        .readdata
		.FFT_STadapter_0_s0_writedata                  (mm_interconnect_0_fft_stadapter_0_s0_writedata),                //                                        .writedata
		.sgdma_from_fft_csr_address                    (mm_interconnect_0_sgdma_from_fft_csr_address),                  //                      sgdma_from_fft_csr.address
		.sgdma_from_fft_csr_write                      (mm_interconnect_0_sgdma_from_fft_csr_write),                    //                                        .write
		.sgdma_from_fft_csr_read                       (mm_interconnect_0_sgdma_from_fft_csr_read),                     //                                        .read
		.sgdma_from_fft_csr_readdata                   (mm_interconnect_0_sgdma_from_fft_csr_readdata),                 //                                        .readdata
		.sgdma_from_fft_csr_writedata                  (mm_interconnect_0_sgdma_from_fft_csr_writedata),                //                                        .writedata
		.sgdma_from_fft_csr_byteenable                 (mm_interconnect_0_sgdma_from_fft_csr_byteenable),               //                                        .byteenable
		.sgdma_from_fft_descriptor_slave_write         (mm_interconnect_0_sgdma_from_fft_descriptor_slave_write),       //         sgdma_from_fft_descriptor_slave.write
		.sgdma_from_fft_descriptor_slave_writedata     (mm_interconnect_0_sgdma_from_fft_descriptor_slave_writedata),   //                                        .writedata
		.sgdma_from_fft_descriptor_slave_byteenable    (mm_interconnect_0_sgdma_from_fft_descriptor_slave_byteenable),  //                                        .byteenable
		.sgdma_from_fft_descriptor_slave_waitrequest   (mm_interconnect_0_sgdma_from_fft_descriptor_slave_waitrequest), //                                        .waitrequest
		.sgdma_from_ram_csr_address                    (mm_interconnect_0_sgdma_from_ram_csr_address),                  //                      sgdma_from_ram_csr.address
		.sgdma_from_ram_csr_write                      (mm_interconnect_0_sgdma_from_ram_csr_write),                    //                                        .write
		.sgdma_from_ram_csr_read                       (mm_interconnect_0_sgdma_from_ram_csr_read),                     //                                        .read
		.sgdma_from_ram_csr_readdata                   (mm_interconnect_0_sgdma_from_ram_csr_readdata),                 //                                        .readdata
		.sgdma_from_ram_csr_writedata                  (mm_interconnect_0_sgdma_from_ram_csr_writedata),                //                                        .writedata
		.sgdma_from_ram_csr_byteenable                 (mm_interconnect_0_sgdma_from_ram_csr_byteenable),               //                                        .byteenable
		.sgdma_from_ram_descriptor_slave_write         (mm_interconnect_0_sgdma_from_ram_descriptor_slave_write),       //         sgdma_from_ram_descriptor_slave.write
		.sgdma_from_ram_descriptor_slave_writedata     (mm_interconnect_0_sgdma_from_ram_descriptor_slave_writedata),   //                                        .writedata
		.sgdma_from_ram_descriptor_slave_byteenable    (mm_interconnect_0_sgdma_from_ram_descriptor_slave_byteenable),  //                                        .byteenable
		.sgdma_from_ram_descriptor_slave_waitrequest   (mm_interconnect_0_sgdma_from_ram_descriptor_slave_waitrequest), //                                        .waitrequest
		.sgdma_to_fft_csr_address                      (mm_interconnect_0_sgdma_to_fft_csr_address),                    //                        sgdma_to_fft_csr.address
		.sgdma_to_fft_csr_write                        (mm_interconnect_0_sgdma_to_fft_csr_write),                      //                                        .write
		.sgdma_to_fft_csr_read                         (mm_interconnect_0_sgdma_to_fft_csr_read),                       //                                        .read
		.sgdma_to_fft_csr_readdata                     (mm_interconnect_0_sgdma_to_fft_csr_readdata),                   //                                        .readdata
		.sgdma_to_fft_csr_writedata                    (mm_interconnect_0_sgdma_to_fft_csr_writedata),                  //                                        .writedata
		.sgdma_to_fft_csr_byteenable                   (mm_interconnect_0_sgdma_to_fft_csr_byteenable),                 //                                        .byteenable
		.sgdma_to_fft_descriptor_slave_write           (mm_interconnect_0_sgdma_to_fft_descriptor_slave_write),         //           sgdma_to_fft_descriptor_slave.write
		.sgdma_to_fft_descriptor_slave_writedata       (mm_interconnect_0_sgdma_to_fft_descriptor_slave_writedata),     //                                        .writedata
		.sgdma_to_fft_descriptor_slave_byteenable      (mm_interconnect_0_sgdma_to_fft_descriptor_slave_byteenable),    //                                        .byteenable
		.sgdma_to_fft_descriptor_slave_waitrequest     (mm_interconnect_0_sgdma_to_fft_descriptor_slave_waitrequest)    //                                        .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign fft_ii_0_source_data = { fft_ii_0_source_real[23:0], fft_ii_0_source_imag[23:0], fft_ii_0_fftpts_out[13:0] };

endmodule
